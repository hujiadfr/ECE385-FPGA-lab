module Bus
(
    input logic GateMARMUX
)