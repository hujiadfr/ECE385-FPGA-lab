module datapath (
    input

    output
)



endmodule