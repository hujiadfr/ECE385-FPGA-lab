// final_soc.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module final_soc (
		output wire [9:0]    bullet_1_x_0_export,    //    bullet_1_x_0.export
		output wire [9:0]    bullet_1_x_1_export,    //    bullet_1_x_1.export
		output wire [9:0]    bullet_1_x_2_export,    //    bullet_1_x_2.export
		output wire [9:0]    bullet_1_x_3_export,    //    bullet_1_x_3.export
		output wire [9:0]    bullet_1_x_4_export,    //    bullet_1_x_4.export
		output wire [9:0]    bullet_1_x_5_export,    //    bullet_1_x_5.export
		output wire [9:0]    bullet_1_x_6_export,    //    bullet_1_x_6.export
		output wire [9:0]    bullet_1_x_7_export,    //    bullet_1_x_7.export
		output wire [9:0]    bullet_1_x_8_export,    //    bullet_1_x_8.export
		output wire [9:0]    bullet_1_x_9_export,    //    bullet_1_x_9.export
		output wire [9:0]    bullet_1_y_0_export,    //    bullet_1_y_0.export
		output wire [9:0]    bullet_1_y_1_export,    //    bullet_1_y_1.export
		output wire [9:0]    bullet_1_y_2_export,    //    bullet_1_y_2.export
		output wire [9:0]    bullet_1_y_3_export,    //    bullet_1_y_3.export
		output wire [9:0]    bullet_1_y_4_export,    //    bullet_1_y_4.export
		output wire [9:0]    bullet_1_y_5_export,    //    bullet_1_y_5.export
		output wire [9:0]    bullet_1_y_6_export,    //    bullet_1_y_6.export
		output wire [9:0]    bullet_1_y_7_export,    //    bullet_1_y_7.export
		output wire [9:0]    bullet_1_y_8_export,    //    bullet_1_y_8.export
		output wire [9:0]    bullet_1_y_9_export,    //    bullet_1_y_9.export
		output wire [9:0]    bullet_2_x_0_export,    //    bullet_2_x_0.export
		output wire [9:0]    bullet_2_x_1_export,    //    bullet_2_x_1.export
		output wire [9:0]    bullet_2_x_2_export,    //    bullet_2_x_2.export
		output wire [9:0]    bullet_2_x_3_export,    //    bullet_2_x_3.export
		output wire [9:0]    bullet_2_x_4_export,    //    bullet_2_x_4.export
		output wire [9:0]    bullet_2_x_5_export,    //    bullet_2_x_5.export
		output wire [9:0]    bullet_2_x_6_export,    //    bullet_2_x_6.export
		output wire [9:0]    bullet_2_x_7_export,    //    bullet_2_x_7.export
		output wire [9:0]    bullet_2_x_8_export,    //    bullet_2_x_8.export
		output wire [9:0]    bullet_2_x_9_export,    //    bullet_2_x_9.export
		output wire [9:0]    bullet_2_y_0_export,    //    bullet_2_y_0.export
		output wire [9:0]    bullet_2_y_1_export,    //    bullet_2_y_1.export
		output wire [9:0]    bullet_2_y_2_export,    //    bullet_2_y_2.export
		output wire [9:0]    bullet_2_y_3_export,    //    bullet_2_y_3.export
		output wire [9:0]    bullet_2_y_4_export,    //    bullet_2_y_4.export
		output wire [9:0]    bullet_2_y_5_export,    //    bullet_2_y_5.export
		output wire [9:0]    bullet_2_y_6_export,    //    bullet_2_y_6.export
		output wire [9:0]    bullet_2_y_7_export,    //    bullet_2_y_7.export
		output wire [9:0]    bullet_2_y_8_export,    //    bullet_2_y_8.export
		output wire [9:0]    bullet_2_y_9_export,    //    bullet_2_y_9.export
		input  wire          clk_clk,                //             clk.clk
		output wire [2047:0] game_readdata,          //            game.readdata
		output wire [7:0]    keycode_0_export,       //       keycode_0.export
		output wire [1:0]    otg_hpi_address_export, // otg_hpi_address.export
		output wire          otg_hpi_cs_export,      //      otg_hpi_cs.export
		input  wire [15:0]   otg_hpi_data_in_port,   //    otg_hpi_data.in_port
		output wire [15:0]   otg_hpi_data_out_port,  //                .out_port
		output wire          otg_hpi_r_export,       //       otg_hpi_r.export
		output wire          otg_hpi_reset_export,   //   otg_hpi_reset.export
		output wire          otg_hpi_w_export,       //       otg_hpi_w.export
		input  wire          reset_reset_n,          //           reset.reset_n
		output wire          sdram_clk_clk,          //       sdram_clk.clk
		output wire [12:0]   sdram_wire_addr,        //      sdram_wire.addr
		output wire [1:0]    sdram_wire_ba,          //                .ba
		output wire          sdram_wire_cas_n,       //                .cas_n
		output wire          sdram_wire_cke,         //                .cke
		output wire          sdram_wire_cs_n,        //                .cs_n
		inout  wire [31:0]   sdram_wire_dq,          //                .dq
		output wire [3:0]    sdram_wire_dqm,         //                .dqm
		output wire          sdram_wire_ras_n,       //                .ras_n
		output wire          sdram_wire_we_n         //                .we_n
	);

	wire         sdram_pll_c0_clk;                                            // sdram_pll:c0 -> [SDRAM:clk, mm_interconnect_0:sdram_pll_c0_clk, rst_controller:clk]
	wire  [31:0] nios2_gen2_0_data_master_readdata;                           // mm_interconnect_0:nios2_gen2_0_data_master_readdata -> nios2_gen2_0:d_readdata
	wire         nios2_gen2_0_data_master_waitrequest;                        // mm_interconnect_0:nios2_gen2_0_data_master_waitrequest -> nios2_gen2_0:d_waitrequest
	wire         nios2_gen2_0_data_master_debugaccess;                        // nios2_gen2_0:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:nios2_gen2_0_data_master_debugaccess
	wire  [28:0] nios2_gen2_0_data_master_address;                            // nios2_gen2_0:d_address -> mm_interconnect_0:nios2_gen2_0_data_master_address
	wire   [3:0] nios2_gen2_0_data_master_byteenable;                         // nios2_gen2_0:d_byteenable -> mm_interconnect_0:nios2_gen2_0_data_master_byteenable
	wire         nios2_gen2_0_data_master_read;                               // nios2_gen2_0:d_read -> mm_interconnect_0:nios2_gen2_0_data_master_read
	wire         nios2_gen2_0_data_master_write;                              // nios2_gen2_0:d_write -> mm_interconnect_0:nios2_gen2_0_data_master_write
	wire  [31:0] nios2_gen2_0_data_master_writedata;                          // nios2_gen2_0:d_writedata -> mm_interconnect_0:nios2_gen2_0_data_master_writedata
	wire  [31:0] nios2_gen2_0_instruction_master_readdata;                    // mm_interconnect_0:nios2_gen2_0_instruction_master_readdata -> nios2_gen2_0:i_readdata
	wire         nios2_gen2_0_instruction_master_waitrequest;                 // mm_interconnect_0:nios2_gen2_0_instruction_master_waitrequest -> nios2_gen2_0:i_waitrequest
	wire  [28:0] nios2_gen2_0_instruction_master_address;                     // nios2_gen2_0:i_address -> mm_interconnect_0:nios2_gen2_0_instruction_master_address
	wire         nios2_gen2_0_instruction_master_read;                        // nios2_gen2_0:i_read -> mm_interconnect_0:nios2_gen2_0_instruction_master_read
	wire         mm_interconnect_0_game_core_game_slave_chipselect;           // mm_interconnect_0:game_core_GAME_Slave_chipselect -> game_core:AVL_CS
	wire  [31:0] mm_interconnect_0_game_core_game_slave_readdata;             // game_core:AVL_READDATA -> mm_interconnect_0:game_core_GAME_Slave_readdata
	wire   [5:0] mm_interconnect_0_game_core_game_slave_address;              // mm_interconnect_0:game_core_GAME_Slave_address -> game_core:AVL_ADDR
	wire         mm_interconnect_0_game_core_game_slave_read;                 // mm_interconnect_0:game_core_GAME_Slave_read -> game_core:AVL_READ
	wire   [3:0] mm_interconnect_0_game_core_game_slave_byteenable;           // mm_interconnect_0:game_core_GAME_Slave_byteenable -> game_core:AVL_BYTE_EN
	wire         mm_interconnect_0_game_core_game_slave_write;                // mm_interconnect_0:game_core_GAME_Slave_write -> game_core:AVL_WRITE
	wire  [31:0] mm_interconnect_0_game_core_game_slave_writedata;            // mm_interconnect_0:game_core_GAME_Slave_writedata -> game_core:AVL_WRITEDATA
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect;  // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_chipselect -> jtag_uart_0:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata;    // jtag_uart_0:av_readdata -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest; // jtag_uart_0:av_waitrequest -> mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address;     // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_address -> jtag_uart_0:av_address
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read;        // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_read -> jtag_uart_0:av_read_n
	wire         mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write;       // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_write -> jtag_uart_0:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata;   // mm_interconnect_0:jtag_uart_0_avalon_jtag_slave_writedata -> jtag_uart_0:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_qsys_0_control_slave_readdata;       // sysid_qsys_0:readdata -> mm_interconnect_0:sysid_qsys_0_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_qsys_0_control_slave_address;        // mm_interconnect_0:sysid_qsys_0_control_slave_address -> sysid_qsys_0:address
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata;     // nios2_gen2_0:debug_mem_slave_readdata -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest;  // nios2_gen2_0:debug_mem_slave_waitrequest -> mm_interconnect_0:nios2_gen2_0_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess;  // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_debugaccess -> nios2_gen2_0:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address;      // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_address -> nios2_gen2_0:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read;         // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_read -> nios2_gen2_0:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable;   // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_byteenable -> nios2_gen2_0:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write;        // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_write -> nios2_gen2_0:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata;    // mm_interconnect_0:nios2_gen2_0_debug_mem_slave_writedata -> nios2_gen2_0:debug_mem_slave_writedata
	wire         mm_interconnect_0_otg_hpi_w_s1_chipselect;                   // mm_interconnect_0:otg_hpi_w_s1_chipselect -> otg_hpi_w:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_readdata;                     // otg_hpi_w:readdata -> mm_interconnect_0:otg_hpi_w_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_w_s1_address;                      // mm_interconnect_0:otg_hpi_w_s1_address -> otg_hpi_w:address
	wire         mm_interconnect_0_otg_hpi_w_s1_write;                        // mm_interconnect_0:otg_hpi_w_s1_write -> otg_hpi_w:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_w_s1_writedata;                    // mm_interconnect_0:otg_hpi_w_s1_writedata -> otg_hpi_w:writedata
	wire         mm_interconnect_0_otg_hpi_r_s1_chipselect;                   // mm_interconnect_0:otg_hpi_r_s1_chipselect -> otg_hpi_r:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_readdata;                     // otg_hpi_r:readdata -> mm_interconnect_0:otg_hpi_r_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_r_s1_address;                      // mm_interconnect_0:otg_hpi_r_s1_address -> otg_hpi_r:address
	wire         mm_interconnect_0_otg_hpi_r_s1_write;                        // mm_interconnect_0:otg_hpi_r_s1_write -> otg_hpi_r:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_r_s1_writedata;                    // mm_interconnect_0:otg_hpi_r_s1_writedata -> otg_hpi_r:writedata
	wire         mm_interconnect_0_otg_hpi_data_s1_chipselect;                // mm_interconnect_0:otg_hpi_data_s1_chipselect -> otg_hpi_data:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_readdata;                  // otg_hpi_data:readdata -> mm_interconnect_0:otg_hpi_data_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_data_s1_address;                   // mm_interconnect_0:otg_hpi_data_s1_address -> otg_hpi_data:address
	wire         mm_interconnect_0_otg_hpi_data_s1_write;                     // mm_interconnect_0:otg_hpi_data_s1_write -> otg_hpi_data:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_data_s1_writedata;                 // mm_interconnect_0:otg_hpi_data_s1_writedata -> otg_hpi_data:writedata
	wire         mm_interconnect_0_otg_hpi_address_s1_chipselect;             // mm_interconnect_0:otg_hpi_address_s1_chipselect -> otg_hpi_address:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_readdata;               // otg_hpi_address:readdata -> mm_interconnect_0:otg_hpi_address_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_address_s1_address;                // mm_interconnect_0:otg_hpi_address_s1_address -> otg_hpi_address:address
	wire         mm_interconnect_0_otg_hpi_address_s1_write;                  // mm_interconnect_0:otg_hpi_address_s1_write -> otg_hpi_address:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_address_s1_writedata;              // mm_interconnect_0:otg_hpi_address_s1_writedata -> otg_hpi_address:writedata
	wire         mm_interconnect_0_otg_hpi_cs_s1_chipselect;                  // mm_interconnect_0:otg_hpi_cs_s1_chipselect -> otg_hpi_cs:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_readdata;                    // otg_hpi_cs:readdata -> mm_interconnect_0:otg_hpi_cs_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_cs_s1_address;                     // mm_interconnect_0:otg_hpi_cs_s1_address -> otg_hpi_cs:address
	wire         mm_interconnect_0_otg_hpi_cs_s1_write;                       // mm_interconnect_0:otg_hpi_cs_s1_write -> otg_hpi_cs:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_cs_s1_writedata;                   // mm_interconnect_0:otg_hpi_cs_s1_writedata -> otg_hpi_cs:writedata
	wire         mm_interconnect_0_otg_hpi_reset_s1_chipselect;               // mm_interconnect_0:otg_hpi_reset_s1_chipselect -> otg_hpi_reset:chipselect
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_readdata;                 // otg_hpi_reset:readdata -> mm_interconnect_0:otg_hpi_reset_s1_readdata
	wire   [1:0] mm_interconnect_0_otg_hpi_reset_s1_address;                  // mm_interconnect_0:otg_hpi_reset_s1_address -> otg_hpi_reset:address
	wire         mm_interconnect_0_otg_hpi_reset_s1_write;                    // mm_interconnect_0:otg_hpi_reset_s1_write -> otg_hpi_reset:write_n
	wire  [31:0] mm_interconnect_0_otg_hpi_reset_s1_writedata;                // mm_interconnect_0:otg_hpi_reset_s1_writedata -> otg_hpi_reset:writedata
	wire         mm_interconnect_0_keycode_0_s1_chipselect;                   // mm_interconnect_0:keycode_0_s1_chipselect -> keycode_0:chipselect
	wire  [31:0] mm_interconnect_0_keycode_0_s1_readdata;                     // keycode_0:readdata -> mm_interconnect_0:keycode_0_s1_readdata
	wire   [1:0] mm_interconnect_0_keycode_0_s1_address;                      // mm_interconnect_0:keycode_0_s1_address -> keycode_0:address
	wire         mm_interconnect_0_keycode_0_s1_write;                        // mm_interconnect_0:keycode_0_s1_write -> keycode_0:write_n
	wire  [31:0] mm_interconnect_0_keycode_0_s1_writedata;                    // mm_interconnect_0:keycode_0_s1_writedata -> keycode_0:writedata
	wire         mm_interconnect_0_sdram_s1_chipselect;                       // mm_interconnect_0:SDRAM_s1_chipselect -> SDRAM:az_cs
	wire  [31:0] mm_interconnect_0_sdram_s1_readdata;                         // SDRAM:za_data -> mm_interconnect_0:SDRAM_s1_readdata
	wire         mm_interconnect_0_sdram_s1_waitrequest;                      // SDRAM:za_waitrequest -> mm_interconnect_0:SDRAM_s1_waitrequest
	wire  [24:0] mm_interconnect_0_sdram_s1_address;                          // mm_interconnect_0:SDRAM_s1_address -> SDRAM:az_addr
	wire         mm_interconnect_0_sdram_s1_read;                             // mm_interconnect_0:SDRAM_s1_read -> SDRAM:az_rd_n
	wire   [3:0] mm_interconnect_0_sdram_s1_byteenable;                       // mm_interconnect_0:SDRAM_s1_byteenable -> SDRAM:az_be_n
	wire         mm_interconnect_0_sdram_s1_readdatavalid;                    // SDRAM:za_valid -> mm_interconnect_0:SDRAM_s1_readdatavalid
	wire         mm_interconnect_0_sdram_s1_write;                            // mm_interconnect_0:SDRAM_s1_write -> SDRAM:az_wr_n
	wire  [31:0] mm_interconnect_0_sdram_s1_writedata;                        // mm_interconnect_0:SDRAM_s1_writedata -> SDRAM:az_data
	wire         mm_interconnect_0_bullet_1_x_0_s1_chipselect;                // mm_interconnect_0:bullet_1_x_0_s1_chipselect -> bullet_1_x_0:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_0_s1_readdata;                  // bullet_1_x_0:readdata -> mm_interconnect_0:bullet_1_x_0_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_0_s1_address;                   // mm_interconnect_0:bullet_1_x_0_s1_address -> bullet_1_x_0:address
	wire         mm_interconnect_0_bullet_1_x_0_s1_write;                     // mm_interconnect_0:bullet_1_x_0_s1_write -> bullet_1_x_0:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_0_s1_writedata;                 // mm_interconnect_0:bullet_1_x_0_s1_writedata -> bullet_1_x_0:writedata
	wire         mm_interconnect_0_bullet_1_x_1_s1_chipselect;                // mm_interconnect_0:bullet_1_x_1_s1_chipselect -> bullet_1_x_1:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_1_s1_readdata;                  // bullet_1_x_1:readdata -> mm_interconnect_0:bullet_1_x_1_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_1_s1_address;                   // mm_interconnect_0:bullet_1_x_1_s1_address -> bullet_1_x_1:address
	wire         mm_interconnect_0_bullet_1_x_1_s1_write;                     // mm_interconnect_0:bullet_1_x_1_s1_write -> bullet_1_x_1:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_1_s1_writedata;                 // mm_interconnect_0:bullet_1_x_1_s1_writedata -> bullet_1_x_1:writedata
	wire         mm_interconnect_0_bullet_1_x_2_s1_chipselect;                // mm_interconnect_0:bullet_1_x_2_s1_chipselect -> bullet_1_x_2:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_2_s1_readdata;                  // bullet_1_x_2:readdata -> mm_interconnect_0:bullet_1_x_2_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_2_s1_address;                   // mm_interconnect_0:bullet_1_x_2_s1_address -> bullet_1_x_2:address
	wire         mm_interconnect_0_bullet_1_x_2_s1_write;                     // mm_interconnect_0:bullet_1_x_2_s1_write -> bullet_1_x_2:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_2_s1_writedata;                 // mm_interconnect_0:bullet_1_x_2_s1_writedata -> bullet_1_x_2:writedata
	wire         mm_interconnect_0_bullet_1_x_3_s1_chipselect;                // mm_interconnect_0:bullet_1_x_3_s1_chipselect -> bullet_1_x_3:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_3_s1_readdata;                  // bullet_1_x_3:readdata -> mm_interconnect_0:bullet_1_x_3_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_3_s1_address;                   // mm_interconnect_0:bullet_1_x_3_s1_address -> bullet_1_x_3:address
	wire         mm_interconnect_0_bullet_1_x_3_s1_write;                     // mm_interconnect_0:bullet_1_x_3_s1_write -> bullet_1_x_3:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_3_s1_writedata;                 // mm_interconnect_0:bullet_1_x_3_s1_writedata -> bullet_1_x_3:writedata
	wire         mm_interconnect_0_bullet_1_x_4_s1_chipselect;                // mm_interconnect_0:bullet_1_x_4_s1_chipselect -> bullet_1_x_4:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_4_s1_readdata;                  // bullet_1_x_4:readdata -> mm_interconnect_0:bullet_1_x_4_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_4_s1_address;                   // mm_interconnect_0:bullet_1_x_4_s1_address -> bullet_1_x_4:address
	wire         mm_interconnect_0_bullet_1_x_4_s1_write;                     // mm_interconnect_0:bullet_1_x_4_s1_write -> bullet_1_x_4:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_4_s1_writedata;                 // mm_interconnect_0:bullet_1_x_4_s1_writedata -> bullet_1_x_4:writedata
	wire         mm_interconnect_0_bullet_1_x_5_s1_chipselect;                // mm_interconnect_0:bullet_1_x_5_s1_chipselect -> bullet_1_x_5:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_5_s1_readdata;                  // bullet_1_x_5:readdata -> mm_interconnect_0:bullet_1_x_5_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_5_s1_address;                   // mm_interconnect_0:bullet_1_x_5_s1_address -> bullet_1_x_5:address
	wire         mm_interconnect_0_bullet_1_x_5_s1_write;                     // mm_interconnect_0:bullet_1_x_5_s1_write -> bullet_1_x_5:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_5_s1_writedata;                 // mm_interconnect_0:bullet_1_x_5_s1_writedata -> bullet_1_x_5:writedata
	wire         mm_interconnect_0_bullet_1_x_6_s1_chipselect;                // mm_interconnect_0:bullet_1_x_6_s1_chipselect -> bullet_1_x_6:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_6_s1_readdata;                  // bullet_1_x_6:readdata -> mm_interconnect_0:bullet_1_x_6_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_6_s1_address;                   // mm_interconnect_0:bullet_1_x_6_s1_address -> bullet_1_x_6:address
	wire         mm_interconnect_0_bullet_1_x_6_s1_write;                     // mm_interconnect_0:bullet_1_x_6_s1_write -> bullet_1_x_6:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_6_s1_writedata;                 // mm_interconnect_0:bullet_1_x_6_s1_writedata -> bullet_1_x_6:writedata
	wire         mm_interconnect_0_bullet_1_x_7_s1_chipselect;                // mm_interconnect_0:bullet_1_x_7_s1_chipselect -> bullet_1_x_7:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_7_s1_readdata;                  // bullet_1_x_7:readdata -> mm_interconnect_0:bullet_1_x_7_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_7_s1_address;                   // mm_interconnect_0:bullet_1_x_7_s1_address -> bullet_1_x_7:address
	wire         mm_interconnect_0_bullet_1_x_7_s1_write;                     // mm_interconnect_0:bullet_1_x_7_s1_write -> bullet_1_x_7:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_7_s1_writedata;                 // mm_interconnect_0:bullet_1_x_7_s1_writedata -> bullet_1_x_7:writedata
	wire         mm_interconnect_0_bullet_1_x_8_s1_chipselect;                // mm_interconnect_0:bullet_1_x_8_s1_chipselect -> bullet_1_x_8:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_8_s1_readdata;                  // bullet_1_x_8:readdata -> mm_interconnect_0:bullet_1_x_8_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_8_s1_address;                   // mm_interconnect_0:bullet_1_x_8_s1_address -> bullet_1_x_8:address
	wire         mm_interconnect_0_bullet_1_x_8_s1_write;                     // mm_interconnect_0:bullet_1_x_8_s1_write -> bullet_1_x_8:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_8_s1_writedata;                 // mm_interconnect_0:bullet_1_x_8_s1_writedata -> bullet_1_x_8:writedata
	wire         mm_interconnect_0_bullet_1_x_9_s1_chipselect;                // mm_interconnect_0:bullet_1_x_9_s1_chipselect -> bullet_1_x_9:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_x_9_s1_readdata;                  // bullet_1_x_9:readdata -> mm_interconnect_0:bullet_1_x_9_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_x_9_s1_address;                   // mm_interconnect_0:bullet_1_x_9_s1_address -> bullet_1_x_9:address
	wire         mm_interconnect_0_bullet_1_x_9_s1_write;                     // mm_interconnect_0:bullet_1_x_9_s1_write -> bullet_1_x_9:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_x_9_s1_writedata;                 // mm_interconnect_0:bullet_1_x_9_s1_writedata -> bullet_1_x_9:writedata
	wire         mm_interconnect_0_bullet_1_y_0_s1_chipselect;                // mm_interconnect_0:bullet_1_y_0_s1_chipselect -> bullet_1_y_0:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_0_s1_readdata;                  // bullet_1_y_0:readdata -> mm_interconnect_0:bullet_1_y_0_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_0_s1_address;                   // mm_interconnect_0:bullet_1_y_0_s1_address -> bullet_1_y_0:address
	wire         mm_interconnect_0_bullet_1_y_0_s1_write;                     // mm_interconnect_0:bullet_1_y_0_s1_write -> bullet_1_y_0:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_0_s1_writedata;                 // mm_interconnect_0:bullet_1_y_0_s1_writedata -> bullet_1_y_0:writedata
	wire         mm_interconnect_0_bullet_1_y_1_s1_chipselect;                // mm_interconnect_0:bullet_1_y_1_s1_chipselect -> bullet_1_y_1:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_1_s1_readdata;                  // bullet_1_y_1:readdata -> mm_interconnect_0:bullet_1_y_1_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_1_s1_address;                   // mm_interconnect_0:bullet_1_y_1_s1_address -> bullet_1_y_1:address
	wire         mm_interconnect_0_bullet_1_y_1_s1_write;                     // mm_interconnect_0:bullet_1_y_1_s1_write -> bullet_1_y_1:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_1_s1_writedata;                 // mm_interconnect_0:bullet_1_y_1_s1_writedata -> bullet_1_y_1:writedata
	wire         mm_interconnect_0_bullet_1_y_2_s1_chipselect;                // mm_interconnect_0:bullet_1_y_2_s1_chipselect -> bullet_1_y_2:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_2_s1_readdata;                  // bullet_1_y_2:readdata -> mm_interconnect_0:bullet_1_y_2_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_2_s1_address;                   // mm_interconnect_0:bullet_1_y_2_s1_address -> bullet_1_y_2:address
	wire         mm_interconnect_0_bullet_1_y_2_s1_write;                     // mm_interconnect_0:bullet_1_y_2_s1_write -> bullet_1_y_2:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_2_s1_writedata;                 // mm_interconnect_0:bullet_1_y_2_s1_writedata -> bullet_1_y_2:writedata
	wire         mm_interconnect_0_bullet_1_y_3_s1_chipselect;                // mm_interconnect_0:bullet_1_y_3_s1_chipselect -> bullet_1_y_3:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_3_s1_readdata;                  // bullet_1_y_3:readdata -> mm_interconnect_0:bullet_1_y_3_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_3_s1_address;                   // mm_interconnect_0:bullet_1_y_3_s1_address -> bullet_1_y_3:address
	wire         mm_interconnect_0_bullet_1_y_3_s1_write;                     // mm_interconnect_0:bullet_1_y_3_s1_write -> bullet_1_y_3:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_3_s1_writedata;                 // mm_interconnect_0:bullet_1_y_3_s1_writedata -> bullet_1_y_3:writedata
	wire         mm_interconnect_0_bullet_1_y_4_s1_chipselect;                // mm_interconnect_0:bullet_1_y_4_s1_chipselect -> bullet_1_y_4:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_4_s1_readdata;                  // bullet_1_y_4:readdata -> mm_interconnect_0:bullet_1_y_4_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_4_s1_address;                   // mm_interconnect_0:bullet_1_y_4_s1_address -> bullet_1_y_4:address
	wire         mm_interconnect_0_bullet_1_y_4_s1_write;                     // mm_interconnect_0:bullet_1_y_4_s1_write -> bullet_1_y_4:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_4_s1_writedata;                 // mm_interconnect_0:bullet_1_y_4_s1_writedata -> bullet_1_y_4:writedata
	wire         mm_interconnect_0_bullet_1_y_5_s1_chipselect;                // mm_interconnect_0:bullet_1_y_5_s1_chipselect -> bullet_1_y_5:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_5_s1_readdata;                  // bullet_1_y_5:readdata -> mm_interconnect_0:bullet_1_y_5_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_5_s1_address;                   // mm_interconnect_0:bullet_1_y_5_s1_address -> bullet_1_y_5:address
	wire         mm_interconnect_0_bullet_1_y_5_s1_write;                     // mm_interconnect_0:bullet_1_y_5_s1_write -> bullet_1_y_5:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_5_s1_writedata;                 // mm_interconnect_0:bullet_1_y_5_s1_writedata -> bullet_1_y_5:writedata
	wire         mm_interconnect_0_bullet_1_y_6_s1_chipselect;                // mm_interconnect_0:bullet_1_y_6_s1_chipselect -> bullet_1_y_6:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_6_s1_readdata;                  // bullet_1_y_6:readdata -> mm_interconnect_0:bullet_1_y_6_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_6_s1_address;                   // mm_interconnect_0:bullet_1_y_6_s1_address -> bullet_1_y_6:address
	wire         mm_interconnect_0_bullet_1_y_6_s1_write;                     // mm_interconnect_0:bullet_1_y_6_s1_write -> bullet_1_y_6:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_6_s1_writedata;                 // mm_interconnect_0:bullet_1_y_6_s1_writedata -> bullet_1_y_6:writedata
	wire         mm_interconnect_0_bullet_1_y_7_s1_chipselect;                // mm_interconnect_0:bullet_1_y_7_s1_chipselect -> bullet_1_y_7:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_7_s1_readdata;                  // bullet_1_y_7:readdata -> mm_interconnect_0:bullet_1_y_7_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_7_s1_address;                   // mm_interconnect_0:bullet_1_y_7_s1_address -> bullet_1_y_7:address
	wire         mm_interconnect_0_bullet_1_y_7_s1_write;                     // mm_interconnect_0:bullet_1_y_7_s1_write -> bullet_1_y_7:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_7_s1_writedata;                 // mm_interconnect_0:bullet_1_y_7_s1_writedata -> bullet_1_y_7:writedata
	wire         mm_interconnect_0_bullet_1_y_8_s1_chipselect;                // mm_interconnect_0:bullet_1_y_8_s1_chipselect -> bullet_1_y_8:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_8_s1_readdata;                  // bullet_1_y_8:readdata -> mm_interconnect_0:bullet_1_y_8_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_8_s1_address;                   // mm_interconnect_0:bullet_1_y_8_s1_address -> bullet_1_y_8:address
	wire         mm_interconnect_0_bullet_1_y_8_s1_write;                     // mm_interconnect_0:bullet_1_y_8_s1_write -> bullet_1_y_8:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_8_s1_writedata;                 // mm_interconnect_0:bullet_1_y_8_s1_writedata -> bullet_1_y_8:writedata
	wire         mm_interconnect_0_bullet_1_y_9_s1_chipselect;                // mm_interconnect_0:bullet_1_y_9_s1_chipselect -> bullet_1_y_9:chipselect
	wire  [31:0] mm_interconnect_0_bullet_1_y_9_s1_readdata;                  // bullet_1_y_9:readdata -> mm_interconnect_0:bullet_1_y_9_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_1_y_9_s1_address;                   // mm_interconnect_0:bullet_1_y_9_s1_address -> bullet_1_y_9:address
	wire         mm_interconnect_0_bullet_1_y_9_s1_write;                     // mm_interconnect_0:bullet_1_y_9_s1_write -> bullet_1_y_9:write_n
	wire  [31:0] mm_interconnect_0_bullet_1_y_9_s1_writedata;                 // mm_interconnect_0:bullet_1_y_9_s1_writedata -> bullet_1_y_9:writedata
	wire         mm_interconnect_0_bullet_2_x_0_s1_chipselect;                // mm_interconnect_0:bullet_2_x_0_s1_chipselect -> bullet_2_x_0:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_0_s1_readdata;                  // bullet_2_x_0:readdata -> mm_interconnect_0:bullet_2_x_0_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_0_s1_address;                   // mm_interconnect_0:bullet_2_x_0_s1_address -> bullet_2_x_0:address
	wire         mm_interconnect_0_bullet_2_x_0_s1_write;                     // mm_interconnect_0:bullet_2_x_0_s1_write -> bullet_2_x_0:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_0_s1_writedata;                 // mm_interconnect_0:bullet_2_x_0_s1_writedata -> bullet_2_x_0:writedata
	wire         mm_interconnect_0_bullet_2_x_1_s1_chipselect;                // mm_interconnect_0:bullet_2_x_1_s1_chipselect -> bullet_2_x_1:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_1_s1_readdata;                  // bullet_2_x_1:readdata -> mm_interconnect_0:bullet_2_x_1_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_1_s1_address;                   // mm_interconnect_0:bullet_2_x_1_s1_address -> bullet_2_x_1:address
	wire         mm_interconnect_0_bullet_2_x_1_s1_write;                     // mm_interconnect_0:bullet_2_x_1_s1_write -> bullet_2_x_1:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_1_s1_writedata;                 // mm_interconnect_0:bullet_2_x_1_s1_writedata -> bullet_2_x_1:writedata
	wire         mm_interconnect_0_bullet_2_x_2_s1_chipselect;                // mm_interconnect_0:bullet_2_x_2_s1_chipselect -> bullet_2_x_2:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_2_s1_readdata;                  // bullet_2_x_2:readdata -> mm_interconnect_0:bullet_2_x_2_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_2_s1_address;                   // mm_interconnect_0:bullet_2_x_2_s1_address -> bullet_2_x_2:address
	wire         mm_interconnect_0_bullet_2_x_2_s1_write;                     // mm_interconnect_0:bullet_2_x_2_s1_write -> bullet_2_x_2:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_2_s1_writedata;                 // mm_interconnect_0:bullet_2_x_2_s1_writedata -> bullet_2_x_2:writedata
	wire         mm_interconnect_0_bullet_2_x_3_s1_chipselect;                // mm_interconnect_0:bullet_2_x_3_s1_chipselect -> bullet_2_x_3:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_3_s1_readdata;                  // bullet_2_x_3:readdata -> mm_interconnect_0:bullet_2_x_3_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_3_s1_address;                   // mm_interconnect_0:bullet_2_x_3_s1_address -> bullet_2_x_3:address
	wire         mm_interconnect_0_bullet_2_x_3_s1_write;                     // mm_interconnect_0:bullet_2_x_3_s1_write -> bullet_2_x_3:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_3_s1_writedata;                 // mm_interconnect_0:bullet_2_x_3_s1_writedata -> bullet_2_x_3:writedata
	wire         mm_interconnect_0_bullet_2_x_4_s1_chipselect;                // mm_interconnect_0:bullet_2_x_4_s1_chipselect -> bullet_2_x_4:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_4_s1_readdata;                  // bullet_2_x_4:readdata -> mm_interconnect_0:bullet_2_x_4_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_4_s1_address;                   // mm_interconnect_0:bullet_2_x_4_s1_address -> bullet_2_x_4:address
	wire         mm_interconnect_0_bullet_2_x_4_s1_write;                     // mm_interconnect_0:bullet_2_x_4_s1_write -> bullet_2_x_4:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_4_s1_writedata;                 // mm_interconnect_0:bullet_2_x_4_s1_writedata -> bullet_2_x_4:writedata
	wire         mm_interconnect_0_bullet_2_x_5_s1_chipselect;                // mm_interconnect_0:bullet_2_x_5_s1_chipselect -> bullet_2_x_5:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_5_s1_readdata;                  // bullet_2_x_5:readdata -> mm_interconnect_0:bullet_2_x_5_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_5_s1_address;                   // mm_interconnect_0:bullet_2_x_5_s1_address -> bullet_2_x_5:address
	wire         mm_interconnect_0_bullet_2_x_5_s1_write;                     // mm_interconnect_0:bullet_2_x_5_s1_write -> bullet_2_x_5:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_5_s1_writedata;                 // mm_interconnect_0:bullet_2_x_5_s1_writedata -> bullet_2_x_5:writedata
	wire         mm_interconnect_0_bullet_2_x_6_s1_chipselect;                // mm_interconnect_0:bullet_2_x_6_s1_chipselect -> bullet_2_x_6:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_6_s1_readdata;                  // bullet_2_x_6:readdata -> mm_interconnect_0:bullet_2_x_6_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_6_s1_address;                   // mm_interconnect_0:bullet_2_x_6_s1_address -> bullet_2_x_6:address
	wire         mm_interconnect_0_bullet_2_x_6_s1_write;                     // mm_interconnect_0:bullet_2_x_6_s1_write -> bullet_2_x_6:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_6_s1_writedata;                 // mm_interconnect_0:bullet_2_x_6_s1_writedata -> bullet_2_x_6:writedata
	wire         mm_interconnect_0_bullet_2_x_7_s1_chipselect;                // mm_interconnect_0:bullet_2_x_7_s1_chipselect -> bullet_2_x_7:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_7_s1_readdata;                  // bullet_2_x_7:readdata -> mm_interconnect_0:bullet_2_x_7_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_7_s1_address;                   // mm_interconnect_0:bullet_2_x_7_s1_address -> bullet_2_x_7:address
	wire         mm_interconnect_0_bullet_2_x_7_s1_write;                     // mm_interconnect_0:bullet_2_x_7_s1_write -> bullet_2_x_7:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_7_s1_writedata;                 // mm_interconnect_0:bullet_2_x_7_s1_writedata -> bullet_2_x_7:writedata
	wire         mm_interconnect_0_bullet_2_x_8_s1_chipselect;                // mm_interconnect_0:bullet_2_x_8_s1_chipselect -> bullet_2_x_8:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_8_s1_readdata;                  // bullet_2_x_8:readdata -> mm_interconnect_0:bullet_2_x_8_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_8_s1_address;                   // mm_interconnect_0:bullet_2_x_8_s1_address -> bullet_2_x_8:address
	wire         mm_interconnect_0_bullet_2_x_8_s1_write;                     // mm_interconnect_0:bullet_2_x_8_s1_write -> bullet_2_x_8:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_8_s1_writedata;                 // mm_interconnect_0:bullet_2_x_8_s1_writedata -> bullet_2_x_8:writedata
	wire         mm_interconnect_0_bullet_2_x_9_s1_chipselect;                // mm_interconnect_0:bullet_2_x_9_s1_chipselect -> bullet_2_x_9:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_x_9_s1_readdata;                  // bullet_2_x_9:readdata -> mm_interconnect_0:bullet_2_x_9_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_x_9_s1_address;                   // mm_interconnect_0:bullet_2_x_9_s1_address -> bullet_2_x_9:address
	wire         mm_interconnect_0_bullet_2_x_9_s1_write;                     // mm_interconnect_0:bullet_2_x_9_s1_write -> bullet_2_x_9:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_x_9_s1_writedata;                 // mm_interconnect_0:bullet_2_x_9_s1_writedata -> bullet_2_x_9:writedata
	wire         mm_interconnect_0_bullet_2_y_0_s1_chipselect;                // mm_interconnect_0:bullet_2_y_0_s1_chipselect -> bullet_2_y_0:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_0_s1_readdata;                  // bullet_2_y_0:readdata -> mm_interconnect_0:bullet_2_y_0_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_0_s1_address;                   // mm_interconnect_0:bullet_2_y_0_s1_address -> bullet_2_y_0:address
	wire         mm_interconnect_0_bullet_2_y_0_s1_write;                     // mm_interconnect_0:bullet_2_y_0_s1_write -> bullet_2_y_0:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_0_s1_writedata;                 // mm_interconnect_0:bullet_2_y_0_s1_writedata -> bullet_2_y_0:writedata
	wire         mm_interconnect_0_bullet_2_y_1_s1_chipselect;                // mm_interconnect_0:bullet_2_y_1_s1_chipselect -> bullet_2_y_1:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_1_s1_readdata;                  // bullet_2_y_1:readdata -> mm_interconnect_0:bullet_2_y_1_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_1_s1_address;                   // mm_interconnect_0:bullet_2_y_1_s1_address -> bullet_2_y_1:address
	wire         mm_interconnect_0_bullet_2_y_1_s1_write;                     // mm_interconnect_0:bullet_2_y_1_s1_write -> bullet_2_y_1:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_1_s1_writedata;                 // mm_interconnect_0:bullet_2_y_1_s1_writedata -> bullet_2_y_1:writedata
	wire         mm_interconnect_0_bullet_2_y_5_s1_chipselect;                // mm_interconnect_0:bullet_2_y_5_s1_chipselect -> bullet_2_y_5:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_5_s1_readdata;                  // bullet_2_y_5:readdata -> mm_interconnect_0:bullet_2_y_5_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_5_s1_address;                   // mm_interconnect_0:bullet_2_y_5_s1_address -> bullet_2_y_5:address
	wire         mm_interconnect_0_bullet_2_y_5_s1_write;                     // mm_interconnect_0:bullet_2_y_5_s1_write -> bullet_2_y_5:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_5_s1_writedata;                 // mm_interconnect_0:bullet_2_y_5_s1_writedata -> bullet_2_y_5:writedata
	wire         mm_interconnect_0_bullet_2_y_6_s1_chipselect;                // mm_interconnect_0:bullet_2_y_6_s1_chipselect -> bullet_2_y_6:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_6_s1_readdata;                  // bullet_2_y_6:readdata -> mm_interconnect_0:bullet_2_y_6_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_6_s1_address;                   // mm_interconnect_0:bullet_2_y_6_s1_address -> bullet_2_y_6:address
	wire         mm_interconnect_0_bullet_2_y_6_s1_write;                     // mm_interconnect_0:bullet_2_y_6_s1_write -> bullet_2_y_6:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_6_s1_writedata;                 // mm_interconnect_0:bullet_2_y_6_s1_writedata -> bullet_2_y_6:writedata
	wire         mm_interconnect_0_bullet_2_y_7_s1_chipselect;                // mm_interconnect_0:bullet_2_y_7_s1_chipselect -> bullet_2_y_7:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_7_s1_readdata;                  // bullet_2_y_7:readdata -> mm_interconnect_0:bullet_2_y_7_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_7_s1_address;                   // mm_interconnect_0:bullet_2_y_7_s1_address -> bullet_2_y_7:address
	wire         mm_interconnect_0_bullet_2_y_7_s1_write;                     // mm_interconnect_0:bullet_2_y_7_s1_write -> bullet_2_y_7:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_7_s1_writedata;                 // mm_interconnect_0:bullet_2_y_7_s1_writedata -> bullet_2_y_7:writedata
	wire         mm_interconnect_0_bullet_2_y_8_s1_chipselect;                // mm_interconnect_0:bullet_2_y_8_s1_chipselect -> bullet_2_y_8:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_8_s1_readdata;                  // bullet_2_y_8:readdata -> mm_interconnect_0:bullet_2_y_8_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_8_s1_address;                   // mm_interconnect_0:bullet_2_y_8_s1_address -> bullet_2_y_8:address
	wire         mm_interconnect_0_bullet_2_y_8_s1_write;                     // mm_interconnect_0:bullet_2_y_8_s1_write -> bullet_2_y_8:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_8_s1_writedata;                 // mm_interconnect_0:bullet_2_y_8_s1_writedata -> bullet_2_y_8:writedata
	wire         mm_interconnect_0_bullet_2_y_9_s1_chipselect;                // mm_interconnect_0:bullet_2_y_9_s1_chipselect -> bullet_2_y_9:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_9_s1_readdata;                  // bullet_2_y_9:readdata -> mm_interconnect_0:bullet_2_y_9_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_9_s1_address;                   // mm_interconnect_0:bullet_2_y_9_s1_address -> bullet_2_y_9:address
	wire         mm_interconnect_0_bullet_2_y_9_s1_write;                     // mm_interconnect_0:bullet_2_y_9_s1_write -> bullet_2_y_9:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_9_s1_writedata;                 // mm_interconnect_0:bullet_2_y_9_s1_writedata -> bullet_2_y_9:writedata
	wire         mm_interconnect_0_bullet_2_y_3_s1_chipselect;                // mm_interconnect_0:bullet_2_y_3_s1_chipselect -> bullet_2_y_3:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_3_s1_readdata;                  // bullet_2_y_3:readdata -> mm_interconnect_0:bullet_2_y_3_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_3_s1_address;                   // mm_interconnect_0:bullet_2_y_3_s1_address -> bullet_2_y_3:address
	wire         mm_interconnect_0_bullet_2_y_3_s1_write;                     // mm_interconnect_0:bullet_2_y_3_s1_write -> bullet_2_y_3:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_3_s1_writedata;                 // mm_interconnect_0:bullet_2_y_3_s1_writedata -> bullet_2_y_3:writedata
	wire         mm_interconnect_0_bullet_2_y_4_s1_chipselect;                // mm_interconnect_0:bullet_2_y_4_s1_chipselect -> bullet_2_y_4:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_4_s1_readdata;                  // bullet_2_y_4:readdata -> mm_interconnect_0:bullet_2_y_4_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_4_s1_address;                   // mm_interconnect_0:bullet_2_y_4_s1_address -> bullet_2_y_4:address
	wire         mm_interconnect_0_bullet_2_y_4_s1_write;                     // mm_interconnect_0:bullet_2_y_4_s1_write -> bullet_2_y_4:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_4_s1_writedata;                 // mm_interconnect_0:bullet_2_y_4_s1_writedata -> bullet_2_y_4:writedata
	wire         mm_interconnect_0_bullet_2_y_2_s1_chipselect;                // mm_interconnect_0:bullet_2_y_2_s1_chipselect -> bullet_2_y_2:chipselect
	wire  [31:0] mm_interconnect_0_bullet_2_y_2_s1_readdata;                  // bullet_2_y_2:readdata -> mm_interconnect_0:bullet_2_y_2_s1_readdata
	wire   [1:0] mm_interconnect_0_bullet_2_y_2_s1_address;                   // mm_interconnect_0:bullet_2_y_2_s1_address -> bullet_2_y_2:address
	wire         mm_interconnect_0_bullet_2_y_2_s1_write;                     // mm_interconnect_0:bullet_2_y_2_s1_write -> bullet_2_y_2:write_n
	wire  [31:0] mm_interconnect_0_bullet_2_y_2_s1_writedata;                 // mm_interconnect_0:bullet_2_y_2_s1_writedata -> bullet_2_y_2:writedata
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_readdata;              // sdram_pll:readdata -> mm_interconnect_0:sdram_pll_pll_slave_readdata
	wire   [1:0] mm_interconnect_0_sdram_pll_pll_slave_address;               // mm_interconnect_0:sdram_pll_pll_slave_address -> sdram_pll:address
	wire         mm_interconnect_0_sdram_pll_pll_slave_read;                  // mm_interconnect_0:sdram_pll_pll_slave_read -> sdram_pll:read
	wire         mm_interconnect_0_sdram_pll_pll_slave_write;                 // mm_interconnect_0:sdram_pll_pll_slave_write -> sdram_pll:write
	wire  [31:0] mm_interconnect_0_sdram_pll_pll_slave_writedata;             // mm_interconnect_0:sdram_pll_pll_slave_writedata -> sdram_pll:writedata
	wire         irq_mapper_receiver0_irq;                                    // jtag_uart_0:av_irq -> irq_mapper:receiver0_irq
	wire  [31:0] nios2_gen2_0_irq_irq;                                        // irq_mapper:sender_irq -> nios2_gen2_0:irq
	wire         rst_controller_reset_out_reset;                              // rst_controller:reset_out -> [SDRAM:reset_n, mm_interconnect_0:SDRAM_reset_reset_bridge_in_reset_reset]
	wire         nios2_gen2_0_debug_reset_request_reset;                      // nios2_gen2_0:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	wire         rst_controller_001_reset_out_reset;                          // rst_controller_001:reset_out -> [bullet_1_x_0:reset_n, bullet_1_x_1:reset_n, bullet_1_x_2:reset_n, bullet_1_x_3:reset_n, bullet_1_x_4:reset_n, bullet_1_x_5:reset_n, bullet_1_x_6:reset_n, bullet_1_x_7:reset_n, bullet_1_x_8:reset_n, bullet_1_x_9:reset_n, bullet_1_y_0:reset_n, bullet_1_y_1:reset_n, bullet_1_y_2:reset_n, bullet_1_y_3:reset_n, bullet_1_y_4:reset_n, bullet_1_y_5:reset_n, bullet_1_y_6:reset_n, bullet_1_y_7:reset_n, bullet_1_y_8:reset_n, bullet_1_y_9:reset_n, bullet_2_x_0:reset_n, bullet_2_x_1:reset_n, bullet_2_x_2:reset_n, bullet_2_x_3:reset_n, bullet_2_x_4:reset_n, bullet_2_x_5:reset_n, bullet_2_x_6:reset_n, bullet_2_x_7:reset_n, bullet_2_x_8:reset_n, bullet_2_x_9:reset_n, bullet_2_y_0:reset_n, bullet_2_y_1:reset_n, bullet_2_y_2:reset_n, bullet_2_y_3:reset_n, bullet_2_y_4:reset_n, bullet_2_y_5:reset_n, bullet_2_y_6:reset_n, bullet_2_y_7:reset_n, bullet_2_y_8:reset_n, bullet_2_y_9:reset_n, game_core:RESET, irq_mapper:reset, jtag_uart_0:rst_n, keycode_0:reset_n, mm_interconnect_0:nios2_gen2_0_reset_reset_bridge_in_reset_reset, nios2_gen2_0:reset_n, otg_hpi_address:reset_n, otg_hpi_cs:reset_n, otg_hpi_data:reset_n, otg_hpi_r:reset_n, otg_hpi_reset:reset_n, otg_hpi_w:reset_n, rst_translator:in_reset, sdram_pll:reset, sysid_qsys_0:reset_n]
	wire         rst_controller_001_reset_out_reset_req;                      // rst_controller_001:reset_req -> [nios2_gen2_0:reset_req, rst_translator:reset_req_in]

	final_soc_SDRAM sdram (
		.clk            (sdram_pll_c0_clk),                         //   clk.clk
		.reset_n        (~rst_controller_reset_out_reset),          // reset.reset_n
		.az_addr        (mm_interconnect_0_sdram_s1_address),       //    s1.address
		.az_be_n        (~mm_interconnect_0_sdram_s1_byteenable),   //      .byteenable_n
		.az_cs          (mm_interconnect_0_sdram_s1_chipselect),    //      .chipselect
		.az_data        (mm_interconnect_0_sdram_s1_writedata),     //      .writedata
		.az_rd_n        (~mm_interconnect_0_sdram_s1_read),         //      .read_n
		.az_wr_n        (~mm_interconnect_0_sdram_s1_write),        //      .write_n
		.za_data        (mm_interconnect_0_sdram_s1_readdata),      //      .readdata
		.za_valid       (mm_interconnect_0_sdram_s1_readdatavalid), //      .readdatavalid
		.za_waitrequest (mm_interconnect_0_sdram_s1_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                          //  wire.export
		.zs_ba          (sdram_wire_ba),                            //      .export
		.zs_cas_n       (sdram_wire_cas_n),                         //      .export
		.zs_cke         (sdram_wire_cke),                           //      .export
		.zs_cs_n        (sdram_wire_cs_n),                          //      .export
		.zs_dq          (sdram_wire_dq),                            //      .export
		.zs_dqm         (sdram_wire_dqm),                           //      .export
		.zs_ras_n       (sdram_wire_ras_n),                         //      .export
		.zs_we_n        (sdram_wire_we_n)                           //      .export
	);

	final_soc_bullet_1_x_0 bullet_1_x_0 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_0_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_0_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_1 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_1_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_1_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_2 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_2_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_2_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_3 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_3_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_3_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_4 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_4_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_4_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_5 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_5_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_5_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_6 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_6_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_6_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_7 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_7_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_7_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_8 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_8_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_8_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_x_9 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_x_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_x_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_x_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_x_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_x_9_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_x_9_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_0 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_0_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_0_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_1 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_1_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_1_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_2 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_2_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_2_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_3 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_3_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_3_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_4 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_4_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_4_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_5 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_5_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_5_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_6 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_6_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_6_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_7 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_7_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_7_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_8 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_8_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_8_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_1_y_9 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_1_y_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_1_y_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_1_y_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_1_y_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_1_y_9_s1_readdata),   //                    .readdata
		.out_port   (bullet_1_y_9_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_0 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_0_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_0_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_1 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_1_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_1_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_2 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_2_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_2_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_3 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_3_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_3_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_4 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_4_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_4_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_5 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_5_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_5_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_6 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_6_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_6_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_7 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_7_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_7_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_8 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_8_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_8_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_x_9 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_x_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_x_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_x_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_x_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_x_9_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_x_9_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_0 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_0_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_0_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_1 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_1_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_1_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_2 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_2_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_2_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_3 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_3_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_3_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_4 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_4_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_4_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_5 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_5_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_5_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_5_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_5_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_5_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_5_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_6 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_6_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_6_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_6_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_6_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_6_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_6_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_7 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_7_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_7_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_7_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_7_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_7_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_7_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_8 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_8_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_8_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_8_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_8_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_8_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_8_export)                           // external_connection.export
	);

	final_soc_bullet_1_x_0 bullet_2_y_9 (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_bullet_2_y_9_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_bullet_2_y_9_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_bullet_2_y_9_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_bullet_2_y_9_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_bullet_2_y_9_s1_readdata),   //                    .readdata
		.out_port   (bullet_2_y_9_export)                           // external_connection.export
	);

	avalon_game_interface game_core (
		.CLK           (clk_clk),                                           //         CLK.clk
		.RESET         (rst_controller_001_reset_out_reset),                //        REST.reset
		.AVL_ADDR      (mm_interconnect_0_game_core_game_slave_address),    //  GAME_Slave.address
		.AVL_BYTE_EN   (mm_interconnect_0_game_core_game_slave_byteenable), //            .byteenable
		.AVL_CS        (mm_interconnect_0_game_core_game_slave_chipselect), //            .chipselect
		.AVL_READ      (mm_interconnect_0_game_core_game_slave_read),       //            .read
		.AVL_READDATA  (mm_interconnect_0_game_core_game_slave_readdata),   //            .readdata
		.AVL_WRITE     (mm_interconnect_0_game_core_game_slave_write),      //            .write
		.AVL_WRITEDATA (mm_interconnect_0_game_core_game_slave_writedata),  //            .writedata
		.EXPORT_DATA   (game_readdata)                                      // conduit_end.readdata
	);

	final_soc_jtag_uart_0 jtag_uart_0 (
		.clk            (clk_clk),                                                     //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                         //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                     //               irq.irq
	);

	final_soc_keycode_0 keycode_0 (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_keycode_0_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_keycode_0_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_keycode_0_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_keycode_0_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_keycode_0_s1_readdata),   //                    .readdata
		.out_port   (keycode_0_export)                           // external_connection.export
	);

	final_soc_nios2_gen2_0 nios2_gen2_0 (
		.clk                                 (clk_clk),                                                    //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),                        //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),                     //                          .reset_req
		.d_address                           (nios2_gen2_0_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_gen2_0_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_gen2_0_data_master_read),                              //                          .read
		.d_readdata                          (nios2_gen2_0_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_gen2_0_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_gen2_0_data_master_write),                             //                          .write
		.d_writedata                         (nios2_gen2_0_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_gen2_0_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_gen2_0_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_gen2_0_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_gen2_0_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_gen2_0_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_gen2_0_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_gen2_0_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                            // custom_instruction_master.readra
	);

	final_soc_otg_hpi_address otg_hpi_address (
		.clk        (clk_clk),                                         //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),             //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_address_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_address_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_address_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_address_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_address_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_address_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_cs (
		.clk        (clk_clk),                                    //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),        //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_cs_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_cs_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_cs_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_cs_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_cs_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_cs_export)                           // external_connection.export
	);

	final_soc_otg_hpi_data otg_hpi_data (
		.clk        (clk_clk),                                      //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),          //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_data_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_data_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_data_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_data_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_data_s1_readdata),   //                    .readdata
		.in_port    (otg_hpi_data_in_port),                         // external_connection.export
		.out_port   (otg_hpi_data_out_port)                         //                    .export
	);

	final_soc_otg_hpi_cs otg_hpi_r (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_r_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_r_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_r_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_r_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_r_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_r_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_reset (
		.clk        (clk_clk),                                       //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),           //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_reset_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_reset_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_reset_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_reset_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_reset_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_reset_export)                           // external_connection.export
	);

	final_soc_otg_hpi_cs otg_hpi_w (
		.clk        (clk_clk),                                   //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),       //               reset.reset_n
		.address    (mm_interconnect_0_otg_hpi_w_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_otg_hpi_w_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_otg_hpi_w_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_otg_hpi_w_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_otg_hpi_w_s1_readdata),   //                    .readdata
		.out_port   (otg_hpi_w_export)                           // external_connection.export
	);

	final_soc_sdram_pll sdram_pll (
		.clk                (clk_clk),                                         //       inclk_interface.clk
		.reset              (rst_controller_001_reset_out_reset),              // inclk_interface_reset.reset
		.read               (mm_interconnect_0_sdram_pll_pll_slave_read),      //             pll_slave.read
		.write              (mm_interconnect_0_sdram_pll_pll_slave_write),     //                      .write
		.address            (mm_interconnect_0_sdram_pll_pll_slave_address),   //                      .address
		.readdata           (mm_interconnect_0_sdram_pll_pll_slave_readdata),  //                      .readdata
		.writedata          (mm_interconnect_0_sdram_pll_pll_slave_writedata), //                      .writedata
		.c0                 (sdram_pll_c0_clk),                                //                    c0.clk
		.c1                 (sdram_clk_clk),                                   //                    c1.clk
		.scandone           (),                                                //           (terminated)
		.scandataout        (),                                                //           (terminated)
		.areset             (1'b0),                                            //           (terminated)
		.locked             (),                                                //           (terminated)
		.phasedone          (),                                                //           (terminated)
		.phasecounterselect (4'b0000),                                         //           (terminated)
		.phaseupdown        (1'b0),                                            //           (terminated)
		.phasestep          (1'b0),                                            //           (terminated)
		.scanclk            (1'b0),                                            //           (terminated)
		.scanclkena         (1'b0),                                            //           (terminated)
		.scandata           (1'b0),                                            //           (terminated)
		.configupdate       (1'b0)                                             //           (terminated)
	);

	final_soc_sysid_qsys_0 sysid_qsys_0 (
		.clock    (clk_clk),                                               //           clk.clk
		.reset_n  (~rst_controller_001_reset_out_reset),                   //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_0_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_0_control_slave_address)   //              .address
	);

	final_soc_mm_interconnect_0 mm_interconnect_0 (
		.clk_0_clk_clk                                  (clk_clk),                                                     //                                clk_0_clk.clk
		.sdram_pll_c0_clk                               (sdram_pll_c0_clk),                                            //                             sdram_pll_c0.clk
		.nios2_gen2_0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                          // nios2_gen2_0_reset_reset_bridge_in_reset.reset
		.SDRAM_reset_reset_bridge_in_reset_reset        (rst_controller_reset_out_reset),                              //        SDRAM_reset_reset_bridge_in_reset.reset
		.nios2_gen2_0_data_master_address               (nios2_gen2_0_data_master_address),                            //                 nios2_gen2_0_data_master.address
		.nios2_gen2_0_data_master_waitrequest           (nios2_gen2_0_data_master_waitrequest),                        //                                         .waitrequest
		.nios2_gen2_0_data_master_byteenable            (nios2_gen2_0_data_master_byteenable),                         //                                         .byteenable
		.nios2_gen2_0_data_master_read                  (nios2_gen2_0_data_master_read),                               //                                         .read
		.nios2_gen2_0_data_master_readdata              (nios2_gen2_0_data_master_readdata),                           //                                         .readdata
		.nios2_gen2_0_data_master_write                 (nios2_gen2_0_data_master_write),                              //                                         .write
		.nios2_gen2_0_data_master_writedata             (nios2_gen2_0_data_master_writedata),                          //                                         .writedata
		.nios2_gen2_0_data_master_debugaccess           (nios2_gen2_0_data_master_debugaccess),                        //                                         .debugaccess
		.nios2_gen2_0_instruction_master_address        (nios2_gen2_0_instruction_master_address),                     //          nios2_gen2_0_instruction_master.address
		.nios2_gen2_0_instruction_master_waitrequest    (nios2_gen2_0_instruction_master_waitrequest),                 //                                         .waitrequest
		.nios2_gen2_0_instruction_master_read           (nios2_gen2_0_instruction_master_read),                        //                                         .read
		.nios2_gen2_0_instruction_master_readdata       (nios2_gen2_0_instruction_master_readdata),                    //                                         .readdata
		.bullet_1_x_0_s1_address                        (mm_interconnect_0_bullet_1_x_0_s1_address),                   //                          bullet_1_x_0_s1.address
		.bullet_1_x_0_s1_write                          (mm_interconnect_0_bullet_1_x_0_s1_write),                     //                                         .write
		.bullet_1_x_0_s1_readdata                       (mm_interconnect_0_bullet_1_x_0_s1_readdata),                  //                                         .readdata
		.bullet_1_x_0_s1_writedata                      (mm_interconnect_0_bullet_1_x_0_s1_writedata),                 //                                         .writedata
		.bullet_1_x_0_s1_chipselect                     (mm_interconnect_0_bullet_1_x_0_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_1_s1_address                        (mm_interconnect_0_bullet_1_x_1_s1_address),                   //                          bullet_1_x_1_s1.address
		.bullet_1_x_1_s1_write                          (mm_interconnect_0_bullet_1_x_1_s1_write),                     //                                         .write
		.bullet_1_x_1_s1_readdata                       (mm_interconnect_0_bullet_1_x_1_s1_readdata),                  //                                         .readdata
		.bullet_1_x_1_s1_writedata                      (mm_interconnect_0_bullet_1_x_1_s1_writedata),                 //                                         .writedata
		.bullet_1_x_1_s1_chipselect                     (mm_interconnect_0_bullet_1_x_1_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_2_s1_address                        (mm_interconnect_0_bullet_1_x_2_s1_address),                   //                          bullet_1_x_2_s1.address
		.bullet_1_x_2_s1_write                          (mm_interconnect_0_bullet_1_x_2_s1_write),                     //                                         .write
		.bullet_1_x_2_s1_readdata                       (mm_interconnect_0_bullet_1_x_2_s1_readdata),                  //                                         .readdata
		.bullet_1_x_2_s1_writedata                      (mm_interconnect_0_bullet_1_x_2_s1_writedata),                 //                                         .writedata
		.bullet_1_x_2_s1_chipselect                     (mm_interconnect_0_bullet_1_x_2_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_3_s1_address                        (mm_interconnect_0_bullet_1_x_3_s1_address),                   //                          bullet_1_x_3_s1.address
		.bullet_1_x_3_s1_write                          (mm_interconnect_0_bullet_1_x_3_s1_write),                     //                                         .write
		.bullet_1_x_3_s1_readdata                       (mm_interconnect_0_bullet_1_x_3_s1_readdata),                  //                                         .readdata
		.bullet_1_x_3_s1_writedata                      (mm_interconnect_0_bullet_1_x_3_s1_writedata),                 //                                         .writedata
		.bullet_1_x_3_s1_chipselect                     (mm_interconnect_0_bullet_1_x_3_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_4_s1_address                        (mm_interconnect_0_bullet_1_x_4_s1_address),                   //                          bullet_1_x_4_s1.address
		.bullet_1_x_4_s1_write                          (mm_interconnect_0_bullet_1_x_4_s1_write),                     //                                         .write
		.bullet_1_x_4_s1_readdata                       (mm_interconnect_0_bullet_1_x_4_s1_readdata),                  //                                         .readdata
		.bullet_1_x_4_s1_writedata                      (mm_interconnect_0_bullet_1_x_4_s1_writedata),                 //                                         .writedata
		.bullet_1_x_4_s1_chipselect                     (mm_interconnect_0_bullet_1_x_4_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_5_s1_address                        (mm_interconnect_0_bullet_1_x_5_s1_address),                   //                          bullet_1_x_5_s1.address
		.bullet_1_x_5_s1_write                          (mm_interconnect_0_bullet_1_x_5_s1_write),                     //                                         .write
		.bullet_1_x_5_s1_readdata                       (mm_interconnect_0_bullet_1_x_5_s1_readdata),                  //                                         .readdata
		.bullet_1_x_5_s1_writedata                      (mm_interconnect_0_bullet_1_x_5_s1_writedata),                 //                                         .writedata
		.bullet_1_x_5_s1_chipselect                     (mm_interconnect_0_bullet_1_x_5_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_6_s1_address                        (mm_interconnect_0_bullet_1_x_6_s1_address),                   //                          bullet_1_x_6_s1.address
		.bullet_1_x_6_s1_write                          (mm_interconnect_0_bullet_1_x_6_s1_write),                     //                                         .write
		.bullet_1_x_6_s1_readdata                       (mm_interconnect_0_bullet_1_x_6_s1_readdata),                  //                                         .readdata
		.bullet_1_x_6_s1_writedata                      (mm_interconnect_0_bullet_1_x_6_s1_writedata),                 //                                         .writedata
		.bullet_1_x_6_s1_chipselect                     (mm_interconnect_0_bullet_1_x_6_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_7_s1_address                        (mm_interconnect_0_bullet_1_x_7_s1_address),                   //                          bullet_1_x_7_s1.address
		.bullet_1_x_7_s1_write                          (mm_interconnect_0_bullet_1_x_7_s1_write),                     //                                         .write
		.bullet_1_x_7_s1_readdata                       (mm_interconnect_0_bullet_1_x_7_s1_readdata),                  //                                         .readdata
		.bullet_1_x_7_s1_writedata                      (mm_interconnect_0_bullet_1_x_7_s1_writedata),                 //                                         .writedata
		.bullet_1_x_7_s1_chipselect                     (mm_interconnect_0_bullet_1_x_7_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_8_s1_address                        (mm_interconnect_0_bullet_1_x_8_s1_address),                   //                          bullet_1_x_8_s1.address
		.bullet_1_x_8_s1_write                          (mm_interconnect_0_bullet_1_x_8_s1_write),                     //                                         .write
		.bullet_1_x_8_s1_readdata                       (mm_interconnect_0_bullet_1_x_8_s1_readdata),                  //                                         .readdata
		.bullet_1_x_8_s1_writedata                      (mm_interconnect_0_bullet_1_x_8_s1_writedata),                 //                                         .writedata
		.bullet_1_x_8_s1_chipselect                     (mm_interconnect_0_bullet_1_x_8_s1_chipselect),                //                                         .chipselect
		.bullet_1_x_9_s1_address                        (mm_interconnect_0_bullet_1_x_9_s1_address),                   //                          bullet_1_x_9_s1.address
		.bullet_1_x_9_s1_write                          (mm_interconnect_0_bullet_1_x_9_s1_write),                     //                                         .write
		.bullet_1_x_9_s1_readdata                       (mm_interconnect_0_bullet_1_x_9_s1_readdata),                  //                                         .readdata
		.bullet_1_x_9_s1_writedata                      (mm_interconnect_0_bullet_1_x_9_s1_writedata),                 //                                         .writedata
		.bullet_1_x_9_s1_chipselect                     (mm_interconnect_0_bullet_1_x_9_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_0_s1_address                        (mm_interconnect_0_bullet_1_y_0_s1_address),                   //                          bullet_1_y_0_s1.address
		.bullet_1_y_0_s1_write                          (mm_interconnect_0_bullet_1_y_0_s1_write),                     //                                         .write
		.bullet_1_y_0_s1_readdata                       (mm_interconnect_0_bullet_1_y_0_s1_readdata),                  //                                         .readdata
		.bullet_1_y_0_s1_writedata                      (mm_interconnect_0_bullet_1_y_0_s1_writedata),                 //                                         .writedata
		.bullet_1_y_0_s1_chipselect                     (mm_interconnect_0_bullet_1_y_0_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_1_s1_address                        (mm_interconnect_0_bullet_1_y_1_s1_address),                   //                          bullet_1_y_1_s1.address
		.bullet_1_y_1_s1_write                          (mm_interconnect_0_bullet_1_y_1_s1_write),                     //                                         .write
		.bullet_1_y_1_s1_readdata                       (mm_interconnect_0_bullet_1_y_1_s1_readdata),                  //                                         .readdata
		.bullet_1_y_1_s1_writedata                      (mm_interconnect_0_bullet_1_y_1_s1_writedata),                 //                                         .writedata
		.bullet_1_y_1_s1_chipselect                     (mm_interconnect_0_bullet_1_y_1_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_2_s1_address                        (mm_interconnect_0_bullet_1_y_2_s1_address),                   //                          bullet_1_y_2_s1.address
		.bullet_1_y_2_s1_write                          (mm_interconnect_0_bullet_1_y_2_s1_write),                     //                                         .write
		.bullet_1_y_2_s1_readdata                       (mm_interconnect_0_bullet_1_y_2_s1_readdata),                  //                                         .readdata
		.bullet_1_y_2_s1_writedata                      (mm_interconnect_0_bullet_1_y_2_s1_writedata),                 //                                         .writedata
		.bullet_1_y_2_s1_chipselect                     (mm_interconnect_0_bullet_1_y_2_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_3_s1_address                        (mm_interconnect_0_bullet_1_y_3_s1_address),                   //                          bullet_1_y_3_s1.address
		.bullet_1_y_3_s1_write                          (mm_interconnect_0_bullet_1_y_3_s1_write),                     //                                         .write
		.bullet_1_y_3_s1_readdata                       (mm_interconnect_0_bullet_1_y_3_s1_readdata),                  //                                         .readdata
		.bullet_1_y_3_s1_writedata                      (mm_interconnect_0_bullet_1_y_3_s1_writedata),                 //                                         .writedata
		.bullet_1_y_3_s1_chipselect                     (mm_interconnect_0_bullet_1_y_3_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_4_s1_address                        (mm_interconnect_0_bullet_1_y_4_s1_address),                   //                          bullet_1_y_4_s1.address
		.bullet_1_y_4_s1_write                          (mm_interconnect_0_bullet_1_y_4_s1_write),                     //                                         .write
		.bullet_1_y_4_s1_readdata                       (mm_interconnect_0_bullet_1_y_4_s1_readdata),                  //                                         .readdata
		.bullet_1_y_4_s1_writedata                      (mm_interconnect_0_bullet_1_y_4_s1_writedata),                 //                                         .writedata
		.bullet_1_y_4_s1_chipselect                     (mm_interconnect_0_bullet_1_y_4_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_5_s1_address                        (mm_interconnect_0_bullet_1_y_5_s1_address),                   //                          bullet_1_y_5_s1.address
		.bullet_1_y_5_s1_write                          (mm_interconnect_0_bullet_1_y_5_s1_write),                     //                                         .write
		.bullet_1_y_5_s1_readdata                       (mm_interconnect_0_bullet_1_y_5_s1_readdata),                  //                                         .readdata
		.bullet_1_y_5_s1_writedata                      (mm_interconnect_0_bullet_1_y_5_s1_writedata),                 //                                         .writedata
		.bullet_1_y_5_s1_chipselect                     (mm_interconnect_0_bullet_1_y_5_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_6_s1_address                        (mm_interconnect_0_bullet_1_y_6_s1_address),                   //                          bullet_1_y_6_s1.address
		.bullet_1_y_6_s1_write                          (mm_interconnect_0_bullet_1_y_6_s1_write),                     //                                         .write
		.bullet_1_y_6_s1_readdata                       (mm_interconnect_0_bullet_1_y_6_s1_readdata),                  //                                         .readdata
		.bullet_1_y_6_s1_writedata                      (mm_interconnect_0_bullet_1_y_6_s1_writedata),                 //                                         .writedata
		.bullet_1_y_6_s1_chipselect                     (mm_interconnect_0_bullet_1_y_6_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_7_s1_address                        (mm_interconnect_0_bullet_1_y_7_s1_address),                   //                          bullet_1_y_7_s1.address
		.bullet_1_y_7_s1_write                          (mm_interconnect_0_bullet_1_y_7_s1_write),                     //                                         .write
		.bullet_1_y_7_s1_readdata                       (mm_interconnect_0_bullet_1_y_7_s1_readdata),                  //                                         .readdata
		.bullet_1_y_7_s1_writedata                      (mm_interconnect_0_bullet_1_y_7_s1_writedata),                 //                                         .writedata
		.bullet_1_y_7_s1_chipselect                     (mm_interconnect_0_bullet_1_y_7_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_8_s1_address                        (mm_interconnect_0_bullet_1_y_8_s1_address),                   //                          bullet_1_y_8_s1.address
		.bullet_1_y_8_s1_write                          (mm_interconnect_0_bullet_1_y_8_s1_write),                     //                                         .write
		.bullet_1_y_8_s1_readdata                       (mm_interconnect_0_bullet_1_y_8_s1_readdata),                  //                                         .readdata
		.bullet_1_y_8_s1_writedata                      (mm_interconnect_0_bullet_1_y_8_s1_writedata),                 //                                         .writedata
		.bullet_1_y_8_s1_chipselect                     (mm_interconnect_0_bullet_1_y_8_s1_chipselect),                //                                         .chipselect
		.bullet_1_y_9_s1_address                        (mm_interconnect_0_bullet_1_y_9_s1_address),                   //                          bullet_1_y_9_s1.address
		.bullet_1_y_9_s1_write                          (mm_interconnect_0_bullet_1_y_9_s1_write),                     //                                         .write
		.bullet_1_y_9_s1_readdata                       (mm_interconnect_0_bullet_1_y_9_s1_readdata),                  //                                         .readdata
		.bullet_1_y_9_s1_writedata                      (mm_interconnect_0_bullet_1_y_9_s1_writedata),                 //                                         .writedata
		.bullet_1_y_9_s1_chipselect                     (mm_interconnect_0_bullet_1_y_9_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_0_s1_address                        (mm_interconnect_0_bullet_2_x_0_s1_address),                   //                          bullet_2_x_0_s1.address
		.bullet_2_x_0_s1_write                          (mm_interconnect_0_bullet_2_x_0_s1_write),                     //                                         .write
		.bullet_2_x_0_s1_readdata                       (mm_interconnect_0_bullet_2_x_0_s1_readdata),                  //                                         .readdata
		.bullet_2_x_0_s1_writedata                      (mm_interconnect_0_bullet_2_x_0_s1_writedata),                 //                                         .writedata
		.bullet_2_x_0_s1_chipselect                     (mm_interconnect_0_bullet_2_x_0_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_1_s1_address                        (mm_interconnect_0_bullet_2_x_1_s1_address),                   //                          bullet_2_x_1_s1.address
		.bullet_2_x_1_s1_write                          (mm_interconnect_0_bullet_2_x_1_s1_write),                     //                                         .write
		.bullet_2_x_1_s1_readdata                       (mm_interconnect_0_bullet_2_x_1_s1_readdata),                  //                                         .readdata
		.bullet_2_x_1_s1_writedata                      (mm_interconnect_0_bullet_2_x_1_s1_writedata),                 //                                         .writedata
		.bullet_2_x_1_s1_chipselect                     (mm_interconnect_0_bullet_2_x_1_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_2_s1_address                        (mm_interconnect_0_bullet_2_x_2_s1_address),                   //                          bullet_2_x_2_s1.address
		.bullet_2_x_2_s1_write                          (mm_interconnect_0_bullet_2_x_2_s1_write),                     //                                         .write
		.bullet_2_x_2_s1_readdata                       (mm_interconnect_0_bullet_2_x_2_s1_readdata),                  //                                         .readdata
		.bullet_2_x_2_s1_writedata                      (mm_interconnect_0_bullet_2_x_2_s1_writedata),                 //                                         .writedata
		.bullet_2_x_2_s1_chipselect                     (mm_interconnect_0_bullet_2_x_2_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_3_s1_address                        (mm_interconnect_0_bullet_2_x_3_s1_address),                   //                          bullet_2_x_3_s1.address
		.bullet_2_x_3_s1_write                          (mm_interconnect_0_bullet_2_x_3_s1_write),                     //                                         .write
		.bullet_2_x_3_s1_readdata                       (mm_interconnect_0_bullet_2_x_3_s1_readdata),                  //                                         .readdata
		.bullet_2_x_3_s1_writedata                      (mm_interconnect_0_bullet_2_x_3_s1_writedata),                 //                                         .writedata
		.bullet_2_x_3_s1_chipselect                     (mm_interconnect_0_bullet_2_x_3_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_4_s1_address                        (mm_interconnect_0_bullet_2_x_4_s1_address),                   //                          bullet_2_x_4_s1.address
		.bullet_2_x_4_s1_write                          (mm_interconnect_0_bullet_2_x_4_s1_write),                     //                                         .write
		.bullet_2_x_4_s1_readdata                       (mm_interconnect_0_bullet_2_x_4_s1_readdata),                  //                                         .readdata
		.bullet_2_x_4_s1_writedata                      (mm_interconnect_0_bullet_2_x_4_s1_writedata),                 //                                         .writedata
		.bullet_2_x_4_s1_chipselect                     (mm_interconnect_0_bullet_2_x_4_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_5_s1_address                        (mm_interconnect_0_bullet_2_x_5_s1_address),                   //                          bullet_2_x_5_s1.address
		.bullet_2_x_5_s1_write                          (mm_interconnect_0_bullet_2_x_5_s1_write),                     //                                         .write
		.bullet_2_x_5_s1_readdata                       (mm_interconnect_0_bullet_2_x_5_s1_readdata),                  //                                         .readdata
		.bullet_2_x_5_s1_writedata                      (mm_interconnect_0_bullet_2_x_5_s1_writedata),                 //                                         .writedata
		.bullet_2_x_5_s1_chipselect                     (mm_interconnect_0_bullet_2_x_5_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_6_s1_address                        (mm_interconnect_0_bullet_2_x_6_s1_address),                   //                          bullet_2_x_6_s1.address
		.bullet_2_x_6_s1_write                          (mm_interconnect_0_bullet_2_x_6_s1_write),                     //                                         .write
		.bullet_2_x_6_s1_readdata                       (mm_interconnect_0_bullet_2_x_6_s1_readdata),                  //                                         .readdata
		.bullet_2_x_6_s1_writedata                      (mm_interconnect_0_bullet_2_x_6_s1_writedata),                 //                                         .writedata
		.bullet_2_x_6_s1_chipselect                     (mm_interconnect_0_bullet_2_x_6_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_7_s1_address                        (mm_interconnect_0_bullet_2_x_7_s1_address),                   //                          bullet_2_x_7_s1.address
		.bullet_2_x_7_s1_write                          (mm_interconnect_0_bullet_2_x_7_s1_write),                     //                                         .write
		.bullet_2_x_7_s1_readdata                       (mm_interconnect_0_bullet_2_x_7_s1_readdata),                  //                                         .readdata
		.bullet_2_x_7_s1_writedata                      (mm_interconnect_0_bullet_2_x_7_s1_writedata),                 //                                         .writedata
		.bullet_2_x_7_s1_chipselect                     (mm_interconnect_0_bullet_2_x_7_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_8_s1_address                        (mm_interconnect_0_bullet_2_x_8_s1_address),                   //                          bullet_2_x_8_s1.address
		.bullet_2_x_8_s1_write                          (mm_interconnect_0_bullet_2_x_8_s1_write),                     //                                         .write
		.bullet_2_x_8_s1_readdata                       (mm_interconnect_0_bullet_2_x_8_s1_readdata),                  //                                         .readdata
		.bullet_2_x_8_s1_writedata                      (mm_interconnect_0_bullet_2_x_8_s1_writedata),                 //                                         .writedata
		.bullet_2_x_8_s1_chipselect                     (mm_interconnect_0_bullet_2_x_8_s1_chipselect),                //                                         .chipselect
		.bullet_2_x_9_s1_address                        (mm_interconnect_0_bullet_2_x_9_s1_address),                   //                          bullet_2_x_9_s1.address
		.bullet_2_x_9_s1_write                          (mm_interconnect_0_bullet_2_x_9_s1_write),                     //                                         .write
		.bullet_2_x_9_s1_readdata                       (mm_interconnect_0_bullet_2_x_9_s1_readdata),                  //                                         .readdata
		.bullet_2_x_9_s1_writedata                      (mm_interconnect_0_bullet_2_x_9_s1_writedata),                 //                                         .writedata
		.bullet_2_x_9_s1_chipselect                     (mm_interconnect_0_bullet_2_x_9_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_0_s1_address                        (mm_interconnect_0_bullet_2_y_0_s1_address),                   //                          bullet_2_y_0_s1.address
		.bullet_2_y_0_s1_write                          (mm_interconnect_0_bullet_2_y_0_s1_write),                     //                                         .write
		.bullet_2_y_0_s1_readdata                       (mm_interconnect_0_bullet_2_y_0_s1_readdata),                  //                                         .readdata
		.bullet_2_y_0_s1_writedata                      (mm_interconnect_0_bullet_2_y_0_s1_writedata),                 //                                         .writedata
		.bullet_2_y_0_s1_chipselect                     (mm_interconnect_0_bullet_2_y_0_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_1_s1_address                        (mm_interconnect_0_bullet_2_y_1_s1_address),                   //                          bullet_2_y_1_s1.address
		.bullet_2_y_1_s1_write                          (mm_interconnect_0_bullet_2_y_1_s1_write),                     //                                         .write
		.bullet_2_y_1_s1_readdata                       (mm_interconnect_0_bullet_2_y_1_s1_readdata),                  //                                         .readdata
		.bullet_2_y_1_s1_writedata                      (mm_interconnect_0_bullet_2_y_1_s1_writedata),                 //                                         .writedata
		.bullet_2_y_1_s1_chipselect                     (mm_interconnect_0_bullet_2_y_1_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_2_s1_address                        (mm_interconnect_0_bullet_2_y_2_s1_address),                   //                          bullet_2_y_2_s1.address
		.bullet_2_y_2_s1_write                          (mm_interconnect_0_bullet_2_y_2_s1_write),                     //                                         .write
		.bullet_2_y_2_s1_readdata                       (mm_interconnect_0_bullet_2_y_2_s1_readdata),                  //                                         .readdata
		.bullet_2_y_2_s1_writedata                      (mm_interconnect_0_bullet_2_y_2_s1_writedata),                 //                                         .writedata
		.bullet_2_y_2_s1_chipselect                     (mm_interconnect_0_bullet_2_y_2_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_3_s1_address                        (mm_interconnect_0_bullet_2_y_3_s1_address),                   //                          bullet_2_y_3_s1.address
		.bullet_2_y_3_s1_write                          (mm_interconnect_0_bullet_2_y_3_s1_write),                     //                                         .write
		.bullet_2_y_3_s1_readdata                       (mm_interconnect_0_bullet_2_y_3_s1_readdata),                  //                                         .readdata
		.bullet_2_y_3_s1_writedata                      (mm_interconnect_0_bullet_2_y_3_s1_writedata),                 //                                         .writedata
		.bullet_2_y_3_s1_chipselect                     (mm_interconnect_0_bullet_2_y_3_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_4_s1_address                        (mm_interconnect_0_bullet_2_y_4_s1_address),                   //                          bullet_2_y_4_s1.address
		.bullet_2_y_4_s1_write                          (mm_interconnect_0_bullet_2_y_4_s1_write),                     //                                         .write
		.bullet_2_y_4_s1_readdata                       (mm_interconnect_0_bullet_2_y_4_s1_readdata),                  //                                         .readdata
		.bullet_2_y_4_s1_writedata                      (mm_interconnect_0_bullet_2_y_4_s1_writedata),                 //                                         .writedata
		.bullet_2_y_4_s1_chipselect                     (mm_interconnect_0_bullet_2_y_4_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_5_s1_address                        (mm_interconnect_0_bullet_2_y_5_s1_address),                   //                          bullet_2_y_5_s1.address
		.bullet_2_y_5_s1_write                          (mm_interconnect_0_bullet_2_y_5_s1_write),                     //                                         .write
		.bullet_2_y_5_s1_readdata                       (mm_interconnect_0_bullet_2_y_5_s1_readdata),                  //                                         .readdata
		.bullet_2_y_5_s1_writedata                      (mm_interconnect_0_bullet_2_y_5_s1_writedata),                 //                                         .writedata
		.bullet_2_y_5_s1_chipselect                     (mm_interconnect_0_bullet_2_y_5_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_6_s1_address                        (mm_interconnect_0_bullet_2_y_6_s1_address),                   //                          bullet_2_y_6_s1.address
		.bullet_2_y_6_s1_write                          (mm_interconnect_0_bullet_2_y_6_s1_write),                     //                                         .write
		.bullet_2_y_6_s1_readdata                       (mm_interconnect_0_bullet_2_y_6_s1_readdata),                  //                                         .readdata
		.bullet_2_y_6_s1_writedata                      (mm_interconnect_0_bullet_2_y_6_s1_writedata),                 //                                         .writedata
		.bullet_2_y_6_s1_chipselect                     (mm_interconnect_0_bullet_2_y_6_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_7_s1_address                        (mm_interconnect_0_bullet_2_y_7_s1_address),                   //                          bullet_2_y_7_s1.address
		.bullet_2_y_7_s1_write                          (mm_interconnect_0_bullet_2_y_7_s1_write),                     //                                         .write
		.bullet_2_y_7_s1_readdata                       (mm_interconnect_0_bullet_2_y_7_s1_readdata),                  //                                         .readdata
		.bullet_2_y_7_s1_writedata                      (mm_interconnect_0_bullet_2_y_7_s1_writedata),                 //                                         .writedata
		.bullet_2_y_7_s1_chipselect                     (mm_interconnect_0_bullet_2_y_7_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_8_s1_address                        (mm_interconnect_0_bullet_2_y_8_s1_address),                   //                          bullet_2_y_8_s1.address
		.bullet_2_y_8_s1_write                          (mm_interconnect_0_bullet_2_y_8_s1_write),                     //                                         .write
		.bullet_2_y_8_s1_readdata                       (mm_interconnect_0_bullet_2_y_8_s1_readdata),                  //                                         .readdata
		.bullet_2_y_8_s1_writedata                      (mm_interconnect_0_bullet_2_y_8_s1_writedata),                 //                                         .writedata
		.bullet_2_y_8_s1_chipselect                     (mm_interconnect_0_bullet_2_y_8_s1_chipselect),                //                                         .chipselect
		.bullet_2_y_9_s1_address                        (mm_interconnect_0_bullet_2_y_9_s1_address),                   //                          bullet_2_y_9_s1.address
		.bullet_2_y_9_s1_write                          (mm_interconnect_0_bullet_2_y_9_s1_write),                     //                                         .write
		.bullet_2_y_9_s1_readdata                       (mm_interconnect_0_bullet_2_y_9_s1_readdata),                  //                                         .readdata
		.bullet_2_y_9_s1_writedata                      (mm_interconnect_0_bullet_2_y_9_s1_writedata),                 //                                         .writedata
		.bullet_2_y_9_s1_chipselect                     (mm_interconnect_0_bullet_2_y_9_s1_chipselect),                //                                         .chipselect
		.game_core_GAME_Slave_address                   (mm_interconnect_0_game_core_game_slave_address),              //                     game_core_GAME_Slave.address
		.game_core_GAME_Slave_write                     (mm_interconnect_0_game_core_game_slave_write),                //                                         .write
		.game_core_GAME_Slave_read                      (mm_interconnect_0_game_core_game_slave_read),                 //                                         .read
		.game_core_GAME_Slave_readdata                  (mm_interconnect_0_game_core_game_slave_readdata),             //                                         .readdata
		.game_core_GAME_Slave_writedata                 (mm_interconnect_0_game_core_game_slave_writedata),            //                                         .writedata
		.game_core_GAME_Slave_byteenable                (mm_interconnect_0_game_core_game_slave_byteenable),           //                                         .byteenable
		.game_core_GAME_Slave_chipselect                (mm_interconnect_0_game_core_game_slave_chipselect),           //                                         .chipselect
		.jtag_uart_0_avalon_jtag_slave_address          (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_address),     //            jtag_uart_0_avalon_jtag_slave.address
		.jtag_uart_0_avalon_jtag_slave_write            (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_write),       //                                         .write
		.jtag_uart_0_avalon_jtag_slave_read             (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_read),        //                                         .read
		.jtag_uart_0_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_readdata),    //                                         .readdata
		.jtag_uart_0_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_writedata),   //                                         .writedata
		.jtag_uart_0_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_waitrequest), //                                         .waitrequest
		.jtag_uart_0_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_uart_0_avalon_jtag_slave_chipselect),  //                                         .chipselect
		.keycode_0_s1_address                           (mm_interconnect_0_keycode_0_s1_address),                      //                             keycode_0_s1.address
		.keycode_0_s1_write                             (mm_interconnect_0_keycode_0_s1_write),                        //                                         .write
		.keycode_0_s1_readdata                          (mm_interconnect_0_keycode_0_s1_readdata),                     //                                         .readdata
		.keycode_0_s1_writedata                         (mm_interconnect_0_keycode_0_s1_writedata),                    //                                         .writedata
		.keycode_0_s1_chipselect                        (mm_interconnect_0_keycode_0_s1_chipselect),                   //                                         .chipselect
		.nios2_gen2_0_debug_mem_slave_address           (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_address),      //             nios2_gen2_0_debug_mem_slave.address
		.nios2_gen2_0_debug_mem_slave_write             (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_write),        //                                         .write
		.nios2_gen2_0_debug_mem_slave_read              (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_read),         //                                         .read
		.nios2_gen2_0_debug_mem_slave_readdata          (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_readdata),     //                                         .readdata
		.nios2_gen2_0_debug_mem_slave_writedata         (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_writedata),    //                                         .writedata
		.nios2_gen2_0_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_byteenable),   //                                         .byteenable
		.nios2_gen2_0_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_waitrequest),  //                                         .waitrequest
		.nios2_gen2_0_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_gen2_0_debug_mem_slave_debugaccess),  //                                         .debugaccess
		.otg_hpi_address_s1_address                     (mm_interconnect_0_otg_hpi_address_s1_address),                //                       otg_hpi_address_s1.address
		.otg_hpi_address_s1_write                       (mm_interconnect_0_otg_hpi_address_s1_write),                  //                                         .write
		.otg_hpi_address_s1_readdata                    (mm_interconnect_0_otg_hpi_address_s1_readdata),               //                                         .readdata
		.otg_hpi_address_s1_writedata                   (mm_interconnect_0_otg_hpi_address_s1_writedata),              //                                         .writedata
		.otg_hpi_address_s1_chipselect                  (mm_interconnect_0_otg_hpi_address_s1_chipselect),             //                                         .chipselect
		.otg_hpi_cs_s1_address                          (mm_interconnect_0_otg_hpi_cs_s1_address),                     //                            otg_hpi_cs_s1.address
		.otg_hpi_cs_s1_write                            (mm_interconnect_0_otg_hpi_cs_s1_write),                       //                                         .write
		.otg_hpi_cs_s1_readdata                         (mm_interconnect_0_otg_hpi_cs_s1_readdata),                    //                                         .readdata
		.otg_hpi_cs_s1_writedata                        (mm_interconnect_0_otg_hpi_cs_s1_writedata),                   //                                         .writedata
		.otg_hpi_cs_s1_chipselect                       (mm_interconnect_0_otg_hpi_cs_s1_chipselect),                  //                                         .chipselect
		.otg_hpi_data_s1_address                        (mm_interconnect_0_otg_hpi_data_s1_address),                   //                          otg_hpi_data_s1.address
		.otg_hpi_data_s1_write                          (mm_interconnect_0_otg_hpi_data_s1_write),                     //                                         .write
		.otg_hpi_data_s1_readdata                       (mm_interconnect_0_otg_hpi_data_s1_readdata),                  //                                         .readdata
		.otg_hpi_data_s1_writedata                      (mm_interconnect_0_otg_hpi_data_s1_writedata),                 //                                         .writedata
		.otg_hpi_data_s1_chipselect                     (mm_interconnect_0_otg_hpi_data_s1_chipselect),                //                                         .chipselect
		.otg_hpi_r_s1_address                           (mm_interconnect_0_otg_hpi_r_s1_address),                      //                             otg_hpi_r_s1.address
		.otg_hpi_r_s1_write                             (mm_interconnect_0_otg_hpi_r_s1_write),                        //                                         .write
		.otg_hpi_r_s1_readdata                          (mm_interconnect_0_otg_hpi_r_s1_readdata),                     //                                         .readdata
		.otg_hpi_r_s1_writedata                         (mm_interconnect_0_otg_hpi_r_s1_writedata),                    //                                         .writedata
		.otg_hpi_r_s1_chipselect                        (mm_interconnect_0_otg_hpi_r_s1_chipselect),                   //                                         .chipselect
		.otg_hpi_reset_s1_address                       (mm_interconnect_0_otg_hpi_reset_s1_address),                  //                         otg_hpi_reset_s1.address
		.otg_hpi_reset_s1_write                         (mm_interconnect_0_otg_hpi_reset_s1_write),                    //                                         .write
		.otg_hpi_reset_s1_readdata                      (mm_interconnect_0_otg_hpi_reset_s1_readdata),                 //                                         .readdata
		.otg_hpi_reset_s1_writedata                     (mm_interconnect_0_otg_hpi_reset_s1_writedata),                //                                         .writedata
		.otg_hpi_reset_s1_chipselect                    (mm_interconnect_0_otg_hpi_reset_s1_chipselect),               //                                         .chipselect
		.otg_hpi_w_s1_address                           (mm_interconnect_0_otg_hpi_w_s1_address),                      //                             otg_hpi_w_s1.address
		.otg_hpi_w_s1_write                             (mm_interconnect_0_otg_hpi_w_s1_write),                        //                                         .write
		.otg_hpi_w_s1_readdata                          (mm_interconnect_0_otg_hpi_w_s1_readdata),                     //                                         .readdata
		.otg_hpi_w_s1_writedata                         (mm_interconnect_0_otg_hpi_w_s1_writedata),                    //                                         .writedata
		.otg_hpi_w_s1_chipselect                        (mm_interconnect_0_otg_hpi_w_s1_chipselect),                   //                                         .chipselect
		.SDRAM_s1_address                               (mm_interconnect_0_sdram_s1_address),                          //                                 SDRAM_s1.address
		.SDRAM_s1_write                                 (mm_interconnect_0_sdram_s1_write),                            //                                         .write
		.SDRAM_s1_read                                  (mm_interconnect_0_sdram_s1_read),                             //                                         .read
		.SDRAM_s1_readdata                              (mm_interconnect_0_sdram_s1_readdata),                         //                                         .readdata
		.SDRAM_s1_writedata                             (mm_interconnect_0_sdram_s1_writedata),                        //                                         .writedata
		.SDRAM_s1_byteenable                            (mm_interconnect_0_sdram_s1_byteenable),                       //                                         .byteenable
		.SDRAM_s1_readdatavalid                         (mm_interconnect_0_sdram_s1_readdatavalid),                    //                                         .readdatavalid
		.SDRAM_s1_waitrequest                           (mm_interconnect_0_sdram_s1_waitrequest),                      //                                         .waitrequest
		.SDRAM_s1_chipselect                            (mm_interconnect_0_sdram_s1_chipselect),                       //                                         .chipselect
		.sdram_pll_pll_slave_address                    (mm_interconnect_0_sdram_pll_pll_slave_address),               //                      sdram_pll_pll_slave.address
		.sdram_pll_pll_slave_write                      (mm_interconnect_0_sdram_pll_pll_slave_write),                 //                                         .write
		.sdram_pll_pll_slave_read                       (mm_interconnect_0_sdram_pll_pll_slave_read),                  //                                         .read
		.sdram_pll_pll_slave_readdata                   (mm_interconnect_0_sdram_pll_pll_slave_readdata),              //                                         .readdata
		.sdram_pll_pll_slave_writedata                  (mm_interconnect_0_sdram_pll_pll_slave_writedata),             //                                         .writedata
		.sysid_qsys_0_control_slave_address             (mm_interconnect_0_sysid_qsys_0_control_slave_address),        //               sysid_qsys_0_control_slave.address
		.sysid_qsys_0_control_slave_readdata            (mm_interconnect_0_sysid_qsys_0_control_slave_readdata)        //                                         .readdata
	);

	final_soc_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.sender_irq    (nios2_gen2_0_irq_irq)                //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (sdram_pll_c0_clk),                       //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),         // reset_out.reset
		.reset_req      (),                                       // (terminated)
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.reset_in1      (nios2_gen2_0_debug_reset_request_reset), // reset_in1.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
