//-------------------------------------------------------------------------
//    Color_Mapper.sv                                                    --
//    Stephen Kempf                                                      --
//    3-1-06                                                             --
//                                                                       --
//    Modified by David Kesler  07-16-2008                               --
//    Translated by Joe Meng    07-07-2013                               --
//    Modified by Po-Han Huang  10-06-2017                               --
//                                                                       --
//    Fall 2017 Distribution                                             --
//                                                                       --
//    For use with ECE 385 Lab 8                                         --
//    University of Illinois ECE Department                              --
//-------------------------------------------------------------------------

// color_mapper: Decide which color to be output to VGA for each pixel.
module  color_mapper ( input              is_ball1, is_ball2,            // Whether current pixel belongs to ball 
                                                              //   or background (computed in ball.sv)
                       input        [11:0] code,
                       input        [9:0] DrawX, DrawY,      // Current pixel coordinates
                       output logic [7:0] VGA_R, VGA_G, VGA_B // VGA RGB output
                     );
    
    logic [7:0] Red, Green, Blue;
    logic [7:0] BRed, BGreen, BBlue;
    logic is_ball;
    palette p(.code(code), .R(BRed), .G(BGreen), .B(BBlue));
    // Output colors to VGA
    logic [7:0] tRed, tGreen, tBlue;
    assign VGA_R = Red;
    assign VGA_G = Green;
    assign VGA_B = Blue;
    
    assign is_ball = is_ball1 || is_ball2;

    // Assign color based on is_ball signal
    always_comb
    begin
        if (is_ball == 1'b1) 
        begin
            // White ball
            Red = 8'hff;
            Green = 8'hff;
            Blue = 8'hff;
        end
        else 
        begin
            // // Background with nice color gradient
            // Red = 8'h3f; 
            // Green = 8'h00;
            // Blue = 8'h7f - {1'b0, DrawX[9:3]};
            Red = BRed;
            Green = BGreen;
            Blue = BBlue;
        end
        //this is for pic background
        
    end 
    
endmodule
