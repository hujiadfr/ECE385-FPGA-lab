module palette (
               input logic [11:0] RGB_12,
               input logic Clk,
               output logic [7:0] R, G, B
               );
					
logic [23:0] out;
assign R = out[23:16];
assign G = out[15:8];
assign B = out[7:0];

always_ff @ (posedge Clk)
    begin
        case (RGB_12)
             12'h000:  out <= 24'h000000;
             12'h001:  out <= 24'h000010;
             12'h002:  out <= 24'h000020;
             12'h003:  out <= 24'h000030;
             12'h004:  out <= 24'h000040;
             12'h005:  out <= 24'h000050;
             12'h006:  out <= 24'h000060;
             12'h007:  out <= 24'h000070;
             12'h008:  out <= 24'h000080;
             12'h009:  out <= 24'h000090;
             12'h00a:  out <= 24'h0000a0;
             12'h00b:  out <= 24'h0000b0;
             12'h00c:  out <= 24'h0000c0;
             12'h00d:  out <= 24'h0000d0;
             12'h00e:  out <= 24'h0000e0;
             12'h00f:  out <= 24'h0000f0;
             12'h010:  out <= 24'h001000;
             12'h011:  out <= 24'h001010;
             12'h012:  out <= 24'h001020;
             12'h013:  out <= 24'h001030;
             12'h014:  out <= 24'h001040;
             12'h015:  out <= 24'h001050;
             12'h016:  out <= 24'h001060;
             12'h017:  out <= 24'h001070;
             12'h018:  out <= 24'h001080;
             12'h019:  out <= 24'h001090;
             12'h01a:  out <= 24'h0010a0;
             12'h01b:  out <= 24'h0010b0;
             12'h01c:  out <= 24'h0010c0;
             12'h01d:  out <= 24'h0010d0;
             12'h01e:  out <= 24'h0010e0;
             12'h01f:  out <= 24'h0010f0;
             12'h020:  out <= 24'h002000;
             12'h021:  out <= 24'h002010;
             12'h022:  out <= 24'h002020;
             12'h023:  out <= 24'h002030;
             12'h024:  out <= 24'h002040;
             12'h025:  out <= 24'h002050;
             12'h026:  out <= 24'h002060;
             12'h027:  out <= 24'h002070;
             12'h028:  out <= 24'h002080;
             12'h029:  out <= 24'h002090;
             12'h02a:  out <= 24'h0020a0;
             12'h02b:  out <= 24'h0020b0;
             12'h02c:  out <= 24'h0020c0;
             12'h02d:  out <= 24'h0020d0;
             12'h02e:  out <= 24'h0020e0;
             12'h02f:  out <= 24'h0020f0;
             12'h030:  out <= 24'h003000;
             12'h031:  out <= 24'h003010;
             12'h032:  out <= 24'h003020;
             12'h033:  out <= 24'h003030;
             12'h034:  out <= 24'h003040;
             12'h035:  out <= 24'h003050;
             12'h036:  out <= 24'h003060;
             12'h037:  out <= 24'h003070;
             12'h038:  out <= 24'h003080;
             12'h039:  out <= 24'h003090;
             12'h03a:  out <= 24'h0030a0;
             12'h03b:  out <= 24'h0030b0;
             12'h03c:  out <= 24'h0030c0;
             12'h03d:  out <= 24'h0030d0;
             12'h03e:  out <= 24'h0030e0;
             12'h03f:  out <= 24'h0030f0;
             12'h040:  out <= 24'h004000;
             12'h041:  out <= 24'h004010;
             12'h042:  out <= 24'h004020;
             12'h043:  out <= 24'h004030;
             12'h044:  out <= 24'h004040;
             12'h045:  out <= 24'h004050;
             12'h046:  out <= 24'h004060;
             12'h047:  out <= 24'h004070;
             12'h048:  out <= 24'h004080;
             12'h049:  out <= 24'h004090;
             12'h04a:  out <= 24'h0040a0;
             12'h04b:  out <= 24'h0040b0;
             12'h04c:  out <= 24'h0040c0;
             12'h04d:  out <= 24'h0040d0;
             12'h04e:  out <= 24'h0040e0;
             12'h04f:  out <= 24'h0040f0;
             12'h050:  out <= 24'h005000;
             12'h051:  out <= 24'h005010;
             12'h052:  out <= 24'h005020;
             12'h053:  out <= 24'h005030;
             12'h054:  out <= 24'h005040;
             12'h055:  out <= 24'h005050;
             12'h056:  out <= 24'h005060;
             12'h057:  out <= 24'h005070;
             12'h058:  out <= 24'h005080;
             12'h059:  out <= 24'h005090;
             12'h05a:  out <= 24'h0050a0;
             12'h05b:  out <= 24'h0050b0;
             12'h05c:  out <= 24'h0050c0;
             12'h05d:  out <= 24'h0050d0;
             12'h05e:  out <= 24'h0050e0;
             12'h05f:  out <= 24'h0050f0;
             12'h060:  out <= 24'h006000;
             12'h061:  out <= 24'h006010;
             12'h062:  out <= 24'h006020;
             12'h063:  out <= 24'h006030;
             12'h064:  out <= 24'h006040;
             12'h065:  out <= 24'h006050;
             12'h066:  out <= 24'h006060;
             12'h067:  out <= 24'h006070;
             12'h068:  out <= 24'h006080;
             12'h069:  out <= 24'h006090;
             12'h06a:  out <= 24'h0060a0;
             12'h06b:  out <= 24'h0060b0;
             12'h06c:  out <= 24'h0060c0;
             12'h06d:  out <= 24'h0060d0;
             12'h06e:  out <= 24'h0060e0;
             12'h06f:  out <= 24'h0060f0;
             12'h070:  out <= 24'h007000;
             12'h071:  out <= 24'h007010;
             12'h072:  out <= 24'h007020;
             12'h073:  out <= 24'h007030;
             12'h074:  out <= 24'h007040;
             12'h075:  out <= 24'h007050;
             12'h076:  out <= 24'h007060;
             12'h077:  out <= 24'h007070;
             12'h078:  out <= 24'h007080;
             12'h079:  out <= 24'h007090;
             12'h07a:  out <= 24'h0070a0;
             12'h07b:  out <= 24'h0070b0;
             12'h07c:  out <= 24'h0070c0;
             12'h07d:  out <= 24'h0070d0;
             12'h07e:  out <= 24'h0070e0;
             12'h07f:  out <= 24'h0070f0;
             12'h080:  out <= 24'h008000;
             12'h081:  out <= 24'h008010;
             12'h082:  out <= 24'h008020;
             12'h083:  out <= 24'h008030;
             12'h084:  out <= 24'h008040;
             12'h085:  out <= 24'h008050;
             12'h086:  out <= 24'h008060;
             12'h087:  out <= 24'h008070;
             12'h088:  out <= 24'h008080;
             12'h089:  out <= 24'h008090;
             12'h08a:  out <= 24'h0080a0;
             12'h08b:  out <= 24'h0080b0;
             12'h08c:  out <= 24'h0080c0;
             12'h08d:  out <= 24'h0080d0;
             12'h08e:  out <= 24'h0080e0;
             12'h08f:  out <= 24'h0080f0;
             12'h090:  out <= 24'h009000;
             12'h091:  out <= 24'h009010;
             12'h092:  out <= 24'h009020;
             12'h093:  out <= 24'h009030;
             12'h094:  out <= 24'h009040;
             12'h095:  out <= 24'h009050;
             12'h096:  out <= 24'h009060;
             12'h097:  out <= 24'h009070;
             12'h098:  out <= 24'h009080;
             12'h099:  out <= 24'h009090;
             12'h09a:  out <= 24'h0090a0;
             12'h09b:  out <= 24'h0090b0;
             12'h09c:  out <= 24'h0090c0;
             12'h09d:  out <= 24'h0090d0;
             12'h09e:  out <= 24'h0090e0;
             12'h09f:  out <= 24'h0090f0;
             12'h0a0:  out <= 24'h00a000;
             12'h0a1:  out <= 24'h00a010;
             12'h0a2:  out <= 24'h00a020;
             12'h0a3:  out <= 24'h00a030;
             12'h0a4:  out <= 24'h00a040;
             12'h0a5:  out <= 24'h00a050;
             12'h0a6:  out <= 24'h00a060;
             12'h0a7:  out <= 24'h00a070;
             12'h0a8:  out <= 24'h00a080;
             12'h0a9:  out <= 24'h00a090;
             12'h0aa:  out <= 24'h00a0a0;
             12'h0ab:  out <= 24'h00a0b0;
             12'h0ac:  out <= 24'h00a0c0;
             12'h0ad:  out <= 24'h00a0d0;
             12'h0ae:  out <= 24'h00a0e0;
             12'h0af:  out <= 24'h00a0f0;
             12'h0b0:  out <= 24'h00b000;
             12'h0b1:  out <= 24'h00b010;
             12'h0b2:  out <= 24'h00b020;
             12'h0b3:  out <= 24'h00b030;
             12'h0b4:  out <= 24'h00b040;
             12'h0b5:  out <= 24'h00b050;
             12'h0b6:  out <= 24'h00b060;
             12'h0b7:  out <= 24'h00b070;
             12'h0b8:  out <= 24'h00b080;
             12'h0b9:  out <= 24'h00b090;
             12'h0ba:  out <= 24'h00b0a0;
             12'h0bb:  out <= 24'h00b0b0;
             12'h0bc:  out <= 24'h00b0c0;
             12'h0bd:  out <= 24'h00b0d0;
             12'h0be:  out <= 24'h00b0e0;
             12'h0bf:  out <= 24'h00b0f0;
             12'h0c0:  out <= 24'h00c000;
             12'h0c1:  out <= 24'h00c010;
             12'h0c2:  out <= 24'h00c020;
             12'h0c3:  out <= 24'h00c030;
             12'h0c4:  out <= 24'h00c040;
             12'h0c5:  out <= 24'h00c050;
             12'h0c6:  out <= 24'h00c060;
             12'h0c7:  out <= 24'h00c070;
             12'h0c8:  out <= 24'h00c080;
             12'h0c9:  out <= 24'h00c090;
             12'h0ca:  out <= 24'h00c0a0;
             12'h0cb:  out <= 24'h00c0b0;
             12'h0cc:  out <= 24'h00c0c0;
             12'h0cd:  out <= 24'h00c0d0;
             12'h0ce:  out <= 24'h00c0e0;
             12'h0cf:  out <= 24'h00c0f0;
             12'h0d0:  out <= 24'h00d000;
             12'h0d1:  out <= 24'h00d010;
             12'h0d2:  out <= 24'h00d020;
             12'h0d3:  out <= 24'h00d030;
             12'h0d4:  out <= 24'h00d040;
             12'h0d5:  out <= 24'h00d050;
             12'h0d6:  out <= 24'h00d060;
             12'h0d7:  out <= 24'h00d070;
             12'h0d8:  out <= 24'h00d080;
             12'h0d9:  out <= 24'h00d090;
             12'h0da:  out <= 24'h00d0a0;
             12'h0db:  out <= 24'h00d0b0;
             12'h0dc:  out <= 24'h00d0c0;
             12'h0dd:  out <= 24'h00d0d0;
             12'h0de:  out <= 24'h00d0e0;
             12'h0df:  out <= 24'h00d0f0;
             12'h0e0:  out <= 24'h00e000;
             12'h0e1:  out <= 24'h00e010;
             12'h0e2:  out <= 24'h00e020;
             12'h0e3:  out <= 24'h00e030;
             12'h0e4:  out <= 24'h00e040;
             12'h0e5:  out <= 24'h00e050;
             12'h0e6:  out <= 24'h00e060;
             12'h0e7:  out <= 24'h00e070;
             12'h0e8:  out <= 24'h00e080;
             12'h0e9:  out <= 24'h00e090;
             12'h0ea:  out <= 24'h00e0a0;
             12'h0eb:  out <= 24'h00e0b0;
             12'h0ec:  out <= 24'h00e0c0;
             12'h0ed:  out <= 24'h00e0d0;
             12'h0ee:  out <= 24'h00e0e0;
             12'h0ef:  out <= 24'h00e0f0;
             12'h0f0:  out <= 24'h00f000;
             12'h0f1:  out <= 24'h00f010;
             12'h0f2:  out <= 24'h00f020;
             12'h0f3:  out <= 24'h00f030;
             12'h0f4:  out <= 24'h00f040;
             12'h0f5:  out <= 24'h00f050;
             12'h0f6:  out <= 24'h00f060;
             12'h0f7:  out <= 24'h00f070;
             12'h0f8:  out <= 24'h00f080;
             12'h0f9:  out <= 24'h00f090;
             12'h0fa:  out <= 24'h00f0a0;
             12'h0fb:  out <= 24'h00f0b0;
             12'h0fc:  out <= 24'h00f0c0;
             12'h0fd:  out <= 24'h00f0d0;
             12'h0fe:  out <= 24'h00f0e0;
             12'h0ff:  out <= 24'h00f0f0;
             12'h100:  out <= 24'h100000;
             12'h101:  out <= 24'h100010;
             12'h102:  out <= 24'h100020;
             12'h103:  out <= 24'h100030;
             12'h104:  out <= 24'h100040;
             12'h105:  out <= 24'h100050;
             12'h106:  out <= 24'h100060;
             12'h107:  out <= 24'h100070;
             12'h108:  out <= 24'h100080;
             12'h109:  out <= 24'h100090;
             12'h10a:  out <= 24'h1000a0;
             12'h10b:  out <= 24'h1000b0;
             12'h10c:  out <= 24'h1000c0;
             12'h10d:  out <= 24'h1000d0;
             12'h10e:  out <= 24'h1000e0;
             12'h10f:  out <= 24'h1000f0;
             12'h110:  out <= 24'h101000;
             12'h111:  out <= 24'h101010;
             12'h112:  out <= 24'h101020;
             12'h113:  out <= 24'h101030;
             12'h114:  out <= 24'h101040;
             12'h115:  out <= 24'h101050;
             12'h116:  out <= 24'h101060;
             12'h117:  out <= 24'h101070;
             12'h118:  out <= 24'h101080;
             12'h119:  out <= 24'h101090;
             12'h11a:  out <= 24'h1010a0;
             12'h11b:  out <= 24'h1010b0;
             12'h11c:  out <= 24'h1010c0;
             12'h11d:  out <= 24'h1010d0;
             12'h11e:  out <= 24'h1010e0;
             12'h11f:  out <= 24'h1010f0;
             12'h120:  out <= 24'h102000;
             12'h121:  out <= 24'h102010;
             12'h122:  out <= 24'h102020;
             12'h123:  out <= 24'h102030;
             12'h124:  out <= 24'h102040;
             12'h125:  out <= 24'h102050;
             12'h126:  out <= 24'h102060;
             12'h127:  out <= 24'h102070;
             12'h128:  out <= 24'h102080;
             12'h129:  out <= 24'h102090;
             12'h12a:  out <= 24'h1020a0;
             12'h12b:  out <= 24'h1020b0;
             12'h12c:  out <= 24'h1020c0;
             12'h12d:  out <= 24'h1020d0;
             12'h12e:  out <= 24'h1020e0;
             12'h12f:  out <= 24'h1020f0;
             12'h130:  out <= 24'h103000;
             12'h131:  out <= 24'h103010;
             12'h132:  out <= 24'h103020;
             12'h133:  out <= 24'h103030;
             12'h134:  out <= 24'h103040;
             12'h135:  out <= 24'h103050;
             12'h136:  out <= 24'h103060;
             12'h137:  out <= 24'h103070;
             12'h138:  out <= 24'h103080;
             12'h139:  out <= 24'h103090;
             12'h13a:  out <= 24'h1030a0;
             12'h13b:  out <= 24'h1030b0;
             12'h13c:  out <= 24'h1030c0;
             12'h13d:  out <= 24'h1030d0;
             12'h13e:  out <= 24'h1030e0;
             12'h13f:  out <= 24'h1030f0;
             12'h140:  out <= 24'h104000;
             12'h141:  out <= 24'h104010;
             12'h142:  out <= 24'h104020;
             12'h143:  out <= 24'h104030;
             12'h144:  out <= 24'h104040;
             12'h145:  out <= 24'h104050;
             12'h146:  out <= 24'h104060;
             12'h147:  out <= 24'h104070;
             12'h148:  out <= 24'h104080;
             12'h149:  out <= 24'h104090;
             12'h14a:  out <= 24'h1040a0;
             12'h14b:  out <= 24'h1040b0;
             12'h14c:  out <= 24'h1040c0;
             12'h14d:  out <= 24'h1040d0;
             12'h14e:  out <= 24'h1040e0;
             12'h14f:  out <= 24'h1040f0;
             12'h150:  out <= 24'h105000;
             12'h151:  out <= 24'h105010;
             12'h152:  out <= 24'h105020;
             12'h153:  out <= 24'h105030;
             12'h154:  out <= 24'h105040;
             12'h155:  out <= 24'h105050;
             12'h156:  out <= 24'h105060;
             12'h157:  out <= 24'h105070;
             12'h158:  out <= 24'h105080;
             12'h159:  out <= 24'h105090;
             12'h15a:  out <= 24'h1050a0;
             12'h15b:  out <= 24'h1050b0;
             12'h15c:  out <= 24'h1050c0;
             12'h15d:  out <= 24'h1050d0;
             12'h15e:  out <= 24'h1050e0;
             12'h15f:  out <= 24'h1050f0;
             12'h160:  out <= 24'h106000;
             12'h161:  out <= 24'h106010;
             12'h162:  out <= 24'h106020;
             12'h163:  out <= 24'h106030;
             12'h164:  out <= 24'h106040;
             12'h165:  out <= 24'h106050;
             12'h166:  out <= 24'h106060;
             12'h167:  out <= 24'h106070;
             12'h168:  out <= 24'h106080;
             12'h169:  out <= 24'h106090;
             12'h16a:  out <= 24'h1060a0;
             12'h16b:  out <= 24'h1060b0;
             12'h16c:  out <= 24'h1060c0;
             12'h16d:  out <= 24'h1060d0;
             12'h16e:  out <= 24'h1060e0;
             12'h16f:  out <= 24'h1060f0;
             12'h170:  out <= 24'h107000;
             12'h171:  out <= 24'h107010;
             12'h172:  out <= 24'h107020;
             12'h173:  out <= 24'h107030;
             12'h174:  out <= 24'h107040;
             12'h175:  out <= 24'h107050;
             12'h176:  out <= 24'h107060;
             12'h177:  out <= 24'h107070;
             12'h178:  out <= 24'h107080;
             12'h179:  out <= 24'h107090;
             12'h17a:  out <= 24'h1070a0;
             12'h17b:  out <= 24'h1070b0;
             12'h17c:  out <= 24'h1070c0;
             12'h17d:  out <= 24'h1070d0;
             12'h17e:  out <= 24'h1070e0;
             12'h17f:  out <= 24'h1070f0;
             12'h180:  out <= 24'h108000;
             12'h181:  out <= 24'h108010;
             12'h182:  out <= 24'h108020;
             12'h183:  out <= 24'h108030;
             12'h184:  out <= 24'h108040;
             12'h185:  out <= 24'h108050;
             12'h186:  out <= 24'h108060;
             12'h187:  out <= 24'h108070;
             12'h188:  out <= 24'h108080;
             12'h189:  out <= 24'h108090;
             12'h18a:  out <= 24'h1080a0;
             12'h18b:  out <= 24'h1080b0;
             12'h18c:  out <= 24'h1080c0;
             12'h18d:  out <= 24'h1080d0;
             12'h18e:  out <= 24'h1080e0;
             12'h18f:  out <= 24'h1080f0;
             12'h190:  out <= 24'h109000;
             12'h191:  out <= 24'h109010;
             12'h192:  out <= 24'h109020;
             12'h193:  out <= 24'h109030;
             12'h194:  out <= 24'h109040;
             12'h195:  out <= 24'h109050;
             12'h196:  out <= 24'h109060;
             12'h197:  out <= 24'h109070;
             12'h198:  out <= 24'h109080;
             12'h199:  out <= 24'h109090;
             12'h19a:  out <= 24'h1090a0;
             12'h19b:  out <= 24'h1090b0;
             12'h19c:  out <= 24'h1090c0;
             12'h19d:  out <= 24'h1090d0;
             12'h19e:  out <= 24'h1090e0;
             12'h19f:  out <= 24'h1090f0;
             12'h1a0:  out <= 24'h10a000;
             12'h1a1:  out <= 24'h10a010;
             12'h1a2:  out <= 24'h10a020;
             12'h1a3:  out <= 24'h10a030;
             12'h1a4:  out <= 24'h10a040;
             12'h1a5:  out <= 24'h10a050;
             12'h1a6:  out <= 24'h10a060;
             12'h1a7:  out <= 24'h10a070;
             12'h1a8:  out <= 24'h10a080;
             12'h1a9:  out <= 24'h10a090;
             12'h1aa:  out <= 24'h10a0a0;
             12'h1ab:  out <= 24'h10a0b0;
             12'h1ac:  out <= 24'h10a0c0;
             12'h1ad:  out <= 24'h10a0d0;
             12'h1ae:  out <= 24'h10a0e0;
             12'h1af:  out <= 24'h10a0f0;
             12'h1b0:  out <= 24'h10b000;
             12'h1b1:  out <= 24'h10b010;
             12'h1b2:  out <= 24'h10b020;
             12'h1b3:  out <= 24'h10b030;
             12'h1b4:  out <= 24'h10b040;
             12'h1b5:  out <= 24'h10b050;
             12'h1b6:  out <= 24'h10b060;
             12'h1b7:  out <= 24'h10b070;
             12'h1b8:  out <= 24'h10b080;
             12'h1b9:  out <= 24'h10b090;
             12'h1ba:  out <= 24'h10b0a0;
             12'h1bb:  out <= 24'h10b0b0;
             12'h1bc:  out <= 24'h10b0c0;
             12'h1bd:  out <= 24'h10b0d0;
             12'h1be:  out <= 24'h10b0e0;
             12'h1bf:  out <= 24'h10b0f0;
             12'h1c0:  out <= 24'h10c000;
             12'h1c1:  out <= 24'h10c010;
             12'h1c2:  out <= 24'h10c020;
             12'h1c3:  out <= 24'h10c030;
             12'h1c4:  out <= 24'h10c040;
             12'h1c5:  out <= 24'h10c050;
             12'h1c6:  out <= 24'h10c060;
             12'h1c7:  out <= 24'h10c070;
             12'h1c8:  out <= 24'h10c080;
             12'h1c9:  out <= 24'h10c090;
             12'h1ca:  out <= 24'h10c0a0;
             12'h1cb:  out <= 24'h10c0b0;
             12'h1cc:  out <= 24'h10c0c0;
             12'h1cd:  out <= 24'h10c0d0;
             12'h1ce:  out <= 24'h10c0e0;
             12'h1cf:  out <= 24'h10c0f0;
             12'h1d0:  out <= 24'h10d000;
             12'h1d1:  out <= 24'h10d010;
             12'h1d2:  out <= 24'h10d020;
             12'h1d3:  out <= 24'h10d030;
             12'h1d4:  out <= 24'h10d040;
             12'h1d5:  out <= 24'h10d050;
             12'h1d6:  out <= 24'h10d060;
             12'h1d7:  out <= 24'h10d070;
             12'h1d8:  out <= 24'h10d080;
             12'h1d9:  out <= 24'h10d090;
             12'h1da:  out <= 24'h10d0a0;
             12'h1db:  out <= 24'h10d0b0;
             12'h1dc:  out <= 24'h10d0c0;
             12'h1dd:  out <= 24'h10d0d0;
             12'h1de:  out <= 24'h10d0e0;
             12'h1df:  out <= 24'h10d0f0;
             12'h1e0:  out <= 24'h10e000;
             12'h1e1:  out <= 24'h10e010;
             12'h1e2:  out <= 24'h10e020;
             12'h1e3:  out <= 24'h10e030;
             12'h1e4:  out <= 24'h10e040;
             12'h1e5:  out <= 24'h10e050;
             12'h1e6:  out <= 24'h10e060;
             12'h1e7:  out <= 24'h10e070;
             12'h1e8:  out <= 24'h10e080;
             12'h1e9:  out <= 24'h10e090;
             12'h1ea:  out <= 24'h10e0a0;
             12'h1eb:  out <= 24'h10e0b0;
             12'h1ec:  out <= 24'h10e0c0;
             12'h1ed:  out <= 24'h10e0d0;
             12'h1ee:  out <= 24'h10e0e0;
             12'h1ef:  out <= 24'h10e0f0;
             12'h1f0:  out <= 24'h10f000;
             12'h1f1:  out <= 24'h10f010;
             12'h1f2:  out <= 24'h10f020;
             12'h1f3:  out <= 24'h10f030;
             12'h1f4:  out <= 24'h10f040;
             12'h1f5:  out <= 24'h10f050;
             12'h1f6:  out <= 24'h10f060;
             12'h1f7:  out <= 24'h10f070;
             12'h1f8:  out <= 24'h10f080;
             12'h1f9:  out <= 24'h10f090;
             12'h1fa:  out <= 24'h10f0a0;
             12'h1fb:  out <= 24'h10f0b0;
             12'h1fc:  out <= 24'h10f0c0;
             12'h1fd:  out <= 24'h10f0d0;
             12'h1fe:  out <= 24'h10f0e0;
             12'h1ff:  out <= 24'h10f0f0;
             12'h200:  out <= 24'h200000;
             12'h201:  out <= 24'h200010;
             12'h202:  out <= 24'h200020;
             12'h203:  out <= 24'h200030;
             12'h204:  out <= 24'h200040;
             12'h205:  out <= 24'h200050;
             12'h206:  out <= 24'h200060;
             12'h207:  out <= 24'h200070;
             12'h208:  out <= 24'h200080;
             12'h209:  out <= 24'h200090;
             12'h20a:  out <= 24'h2000a0;
             12'h20b:  out <= 24'h2000b0;
             12'h20c:  out <= 24'h2000c0;
             12'h20d:  out <= 24'h2000d0;
             12'h20e:  out <= 24'h2000e0;
             12'h20f:  out <= 24'h2000f0;
             12'h210:  out <= 24'h201000;
             12'h211:  out <= 24'h201010;
             12'h212:  out <= 24'h201020;
             12'h213:  out <= 24'h201030;
             12'h214:  out <= 24'h201040;
             12'h215:  out <= 24'h201050;
             12'h216:  out <= 24'h201060;
             12'h217:  out <= 24'h201070;
             12'h218:  out <= 24'h201080;
             12'h219:  out <= 24'h201090;
             12'h21a:  out <= 24'h2010a0;
             12'h21b:  out <= 24'h2010b0;
             12'h21c:  out <= 24'h2010c0;
             12'h21d:  out <= 24'h2010d0;
             12'h21e:  out <= 24'h2010e0;
             12'h21f:  out <= 24'h2010f0;
             12'h220:  out <= 24'h202000;
             12'h221:  out <= 24'h202010;
             12'h222:  out <= 24'h202020;
             12'h223:  out <= 24'h202030;
             12'h224:  out <= 24'h202040;
             12'h225:  out <= 24'h202050;
             12'h226:  out <= 24'h202060;
             12'h227:  out <= 24'h202070;
             12'h228:  out <= 24'h202080;
             12'h229:  out <= 24'h202090;
             12'h22a:  out <= 24'h2020a0;
             12'h22b:  out <= 24'h2020b0;
             12'h22c:  out <= 24'h2020c0;
             12'h22d:  out <= 24'h2020d0;
             12'h22e:  out <= 24'h2020e0;
             12'h22f:  out <= 24'h2020f0;
             12'h230:  out <= 24'h203000;
             12'h231:  out <= 24'h203010;
             12'h232:  out <= 24'h203020;
             12'h233:  out <= 24'h203030;
             12'h234:  out <= 24'h203040;
             12'h235:  out <= 24'h203050;
             12'h236:  out <= 24'h203060;
             12'h237:  out <= 24'h203070;
             12'h238:  out <= 24'h203080;
             12'h239:  out <= 24'h203090;
             12'h23a:  out <= 24'h2030a0;
             12'h23b:  out <= 24'h2030b0;
             12'h23c:  out <= 24'h2030c0;
             12'h23d:  out <= 24'h2030d0;
             12'h23e:  out <= 24'h2030e0;
             12'h23f:  out <= 24'h2030f0;
             12'h240:  out <= 24'h204000;
             12'h241:  out <= 24'h204010;
             12'h242:  out <= 24'h204020;
             12'h243:  out <= 24'h204030;
             12'h244:  out <= 24'h204040;
             12'h245:  out <= 24'h204050;
             12'h246:  out <= 24'h204060;
             12'h247:  out <= 24'h204070;
             12'h248:  out <= 24'h204080;
             12'h249:  out <= 24'h204090;
             12'h24a:  out <= 24'h2040a0;
             12'h24b:  out <= 24'h2040b0;
             12'h24c:  out <= 24'h2040c0;
             12'h24d:  out <= 24'h2040d0;
             12'h24e:  out <= 24'h2040e0;
             12'h24f:  out <= 24'h2040f0;
             12'h250:  out <= 24'h205000;
             12'h251:  out <= 24'h205010;
             12'h252:  out <= 24'h205020;
             12'h253:  out <= 24'h205030;
             12'h254:  out <= 24'h205040;
             12'h255:  out <= 24'h205050;
             12'h256:  out <= 24'h205060;
             12'h257:  out <= 24'h205070;
             12'h258:  out <= 24'h205080;
             12'h259:  out <= 24'h205090;
             12'h25a:  out <= 24'h2050a0;
             12'h25b:  out <= 24'h2050b0;
             12'h25c:  out <= 24'h2050c0;
             12'h25d:  out <= 24'h2050d0;
             12'h25e:  out <= 24'h2050e0;
             12'h25f:  out <= 24'h2050f0;
             12'h260:  out <= 24'h206000;
             12'h261:  out <= 24'h206010;
             12'h262:  out <= 24'h206020;
             12'h263:  out <= 24'h206030;
             12'h264:  out <= 24'h206040;
             12'h265:  out <= 24'h206050;
             12'h266:  out <= 24'h206060;
             12'h267:  out <= 24'h206070;
             12'h268:  out <= 24'h206080;
             12'h269:  out <= 24'h206090;
             12'h26a:  out <= 24'h2060a0;
             12'h26b:  out <= 24'h2060b0;
             12'h26c:  out <= 24'h2060c0;
             12'h26d:  out <= 24'h2060d0;
             12'h26e:  out <= 24'h2060e0;
             12'h26f:  out <= 24'h2060f0;
             12'h270:  out <= 24'h207000;
             12'h271:  out <= 24'h207010;
             12'h272:  out <= 24'h207020;
             12'h273:  out <= 24'h207030;
             12'h274:  out <= 24'h207040;
             12'h275:  out <= 24'h207050;
             12'h276:  out <= 24'h207060;
             12'h277:  out <= 24'h207070;
             12'h278:  out <= 24'h207080;
             12'h279:  out <= 24'h207090;
             12'h27a:  out <= 24'h2070a0;
             12'h27b:  out <= 24'h2070b0;
             12'h27c:  out <= 24'h2070c0;
             12'h27d:  out <= 24'h2070d0;
             12'h27e:  out <= 24'h2070e0;
             12'h27f:  out <= 24'h2070f0;
             12'h280:  out <= 24'h208000;
             12'h281:  out <= 24'h208010;
             12'h282:  out <= 24'h208020;
             12'h283:  out <= 24'h208030;
             12'h284:  out <= 24'h208040;
             12'h285:  out <= 24'h208050;
             12'h286:  out <= 24'h208060;
             12'h287:  out <= 24'h208070;
             12'h288:  out <= 24'h208080;
             12'h289:  out <= 24'h208090;
             12'h28a:  out <= 24'h2080a0;
             12'h28b:  out <= 24'h2080b0;
             12'h28c:  out <= 24'h2080c0;
             12'h28d:  out <= 24'h2080d0;
             12'h28e:  out <= 24'h2080e0;
             12'h28f:  out <= 24'h2080f0;
             12'h290:  out <= 24'h209000;
             12'h291:  out <= 24'h209010;
             12'h292:  out <= 24'h209020;
             12'h293:  out <= 24'h209030;
             12'h294:  out <= 24'h209040;
             12'h295:  out <= 24'h209050;
             12'h296:  out <= 24'h209060;
             12'h297:  out <= 24'h209070;
             12'h298:  out <= 24'h209080;
             12'h299:  out <= 24'h209090;
             12'h29a:  out <= 24'h2090a0;
             12'h29b:  out <= 24'h2090b0;
             12'h29c:  out <= 24'h2090c0;
             12'h29d:  out <= 24'h2090d0;
             12'h29e:  out <= 24'h2090e0;
             12'h29f:  out <= 24'h2090f0;
             12'h2a0:  out <= 24'h20a000;
             12'h2a1:  out <= 24'h20a010;
             12'h2a2:  out <= 24'h20a020;
             12'h2a3:  out <= 24'h20a030;
             12'h2a4:  out <= 24'h20a040;
             12'h2a5:  out <= 24'h20a050;
             12'h2a6:  out <= 24'h20a060;
             12'h2a7:  out <= 24'h20a070;
             12'h2a8:  out <= 24'h20a080;
             12'h2a9:  out <= 24'h20a090;
             12'h2aa:  out <= 24'h20a0a0;
             12'h2ab:  out <= 24'h20a0b0;
             12'h2ac:  out <= 24'h20a0c0;
             12'h2ad:  out <= 24'h20a0d0;
             12'h2ae:  out <= 24'h20a0e0;
             12'h2af:  out <= 24'h20a0f0;
             12'h2b0:  out <= 24'h20b000;
             12'h2b1:  out <= 24'h20b010;
             12'h2b2:  out <= 24'h20b020;
             12'h2b3:  out <= 24'h20b030;
             12'h2b4:  out <= 24'h20b040;
             12'h2b5:  out <= 24'h20b050;
             12'h2b6:  out <= 24'h20b060;
             12'h2b7:  out <= 24'h20b070;
             12'h2b8:  out <= 24'h20b080;
             12'h2b9:  out <= 24'h20b090;
             12'h2ba:  out <= 24'h20b0a0;
             12'h2bb:  out <= 24'h20b0b0;
             12'h2bc:  out <= 24'h20b0c0;
             12'h2bd:  out <= 24'h20b0d0;
             12'h2be:  out <= 24'h20b0e0;
             12'h2bf:  out <= 24'h20b0f0;
             12'h2c0:  out <= 24'h20c000;
             12'h2c1:  out <= 24'h20c010;
             12'h2c2:  out <= 24'h20c020;
             12'h2c3:  out <= 24'h20c030;
             12'h2c4:  out <= 24'h20c040;
             12'h2c5:  out <= 24'h20c050;
             12'h2c6:  out <= 24'h20c060;
             12'h2c7:  out <= 24'h20c070;
             12'h2c8:  out <= 24'h20c080;
             12'h2c9:  out <= 24'h20c090;
             12'h2ca:  out <= 24'h20c0a0;
             12'h2cb:  out <= 24'h20c0b0;
             12'h2cc:  out <= 24'h20c0c0;
             12'h2cd:  out <= 24'h20c0d0;
             12'h2ce:  out <= 24'h20c0e0;
             12'h2cf:  out <= 24'h20c0f0;
             12'h2d0:  out <= 24'h20d000;
             12'h2d1:  out <= 24'h20d010;
             12'h2d2:  out <= 24'h20d020;
             12'h2d3:  out <= 24'h20d030;
             12'h2d4:  out <= 24'h20d040;
             12'h2d5:  out <= 24'h20d050;
             12'h2d6:  out <= 24'h20d060;
             12'h2d7:  out <= 24'h20d070;
             12'h2d8:  out <= 24'h20d080;
             12'h2d9:  out <= 24'h20d090;
             12'h2da:  out <= 24'h20d0a0;
             12'h2db:  out <= 24'h20d0b0;
             12'h2dc:  out <= 24'h20d0c0;
             12'h2dd:  out <= 24'h20d0d0;
             12'h2de:  out <= 24'h20d0e0;
             12'h2df:  out <= 24'h20d0f0;
             12'h2e0:  out <= 24'h20e000;
             12'h2e1:  out <= 24'h20e010;
             12'h2e2:  out <= 24'h20e020;
             12'h2e3:  out <= 24'h20e030;
             12'h2e4:  out <= 24'h20e040;
             12'h2e5:  out <= 24'h20e050;
             12'h2e6:  out <= 24'h20e060;
             12'h2e7:  out <= 24'h20e070;
             12'h2e8:  out <= 24'h20e080;
             12'h2e9:  out <= 24'h20e090;
             12'h2ea:  out <= 24'h20e0a0;
             12'h2eb:  out <= 24'h20e0b0;
             12'h2ec:  out <= 24'h20e0c0;
             12'h2ed:  out <= 24'h20e0d0;
             12'h2ee:  out <= 24'h20e0e0;
             12'h2ef:  out <= 24'h20e0f0;
             12'h2f0:  out <= 24'h20f000;
             12'h2f1:  out <= 24'h20f010;
             12'h2f2:  out <= 24'h20f020;
             12'h2f3:  out <= 24'h20f030;
             12'h2f4:  out <= 24'h20f040;
             12'h2f5:  out <= 24'h20f050;
             12'h2f6:  out <= 24'h20f060;
             12'h2f7:  out <= 24'h20f070;
             12'h2f8:  out <= 24'h20f080;
             12'h2f9:  out <= 24'h20f090;
             12'h2fa:  out <= 24'h20f0a0;
             12'h2fb:  out <= 24'h20f0b0;
             12'h2fc:  out <= 24'h20f0c0;
             12'h2fd:  out <= 24'h20f0d0;
             12'h2fe:  out <= 24'h20f0e0;
             12'h2ff:  out <= 24'h20f0f0;
             12'h300:  out <= 24'h300000;
             12'h301:  out <= 24'h300010;
             12'h302:  out <= 24'h300020;
             12'h303:  out <= 24'h300030;
             12'h304:  out <= 24'h300040;
             12'h305:  out <= 24'h300050;
             12'h306:  out <= 24'h300060;
             12'h307:  out <= 24'h300070;
             12'h308:  out <= 24'h300080;
             12'h309:  out <= 24'h300090;
             12'h30a:  out <= 24'h3000a0;
             12'h30b:  out <= 24'h3000b0;
             12'h30c:  out <= 24'h3000c0;
             12'h30d:  out <= 24'h3000d0;
             12'h30e:  out <= 24'h3000e0;
             12'h30f:  out <= 24'h3000f0;
             12'h310:  out <= 24'h301000;
             12'h311:  out <= 24'h301010;
             12'h312:  out <= 24'h301020;
             12'h313:  out <= 24'h301030;
             12'h314:  out <= 24'h301040;
             12'h315:  out <= 24'h301050;
             12'h316:  out <= 24'h301060;
             12'h317:  out <= 24'h301070;
             12'h318:  out <= 24'h301080;
             12'h319:  out <= 24'h301090;
             12'h31a:  out <= 24'h3010a0;
             12'h31b:  out <= 24'h3010b0;
             12'h31c:  out <= 24'h3010c0;
             12'h31d:  out <= 24'h3010d0;
             12'h31e:  out <= 24'h3010e0;
             12'h31f:  out <= 24'h3010f0;
             12'h320:  out <= 24'h302000;
             12'h321:  out <= 24'h302010;
             12'h322:  out <= 24'h302020;
             12'h323:  out <= 24'h302030;
             12'h324:  out <= 24'h302040;
             12'h325:  out <= 24'h302050;
             12'h326:  out <= 24'h302060;
             12'h327:  out <= 24'h302070;
             12'h328:  out <= 24'h302080;
             12'h329:  out <= 24'h302090;
             12'h32a:  out <= 24'h3020a0;
             12'h32b:  out <= 24'h3020b0;
             12'h32c:  out <= 24'h3020c0;
             12'h32d:  out <= 24'h3020d0;
             12'h32e:  out <= 24'h3020e0;
             12'h32f:  out <= 24'h3020f0;
             12'h330:  out <= 24'h303000;
             12'h331:  out <= 24'h303010;
             12'h332:  out <= 24'h303020;
             12'h333:  out <= 24'h303030;
             12'h334:  out <= 24'h303040;
             12'h335:  out <= 24'h303050;
             12'h336:  out <= 24'h303060;
             12'h337:  out <= 24'h303070;
             12'h338:  out <= 24'h303080;
             12'h339:  out <= 24'h303090;
             12'h33a:  out <= 24'h3030a0;
             12'h33b:  out <= 24'h3030b0;
             12'h33c:  out <= 24'h3030c0;
             12'h33d:  out <= 24'h3030d0;
             12'h33e:  out <= 24'h3030e0;
             12'h33f:  out <= 24'h3030f0;
             12'h340:  out <= 24'h304000;
             12'h341:  out <= 24'h304010;
             12'h342:  out <= 24'h304020;
             12'h343:  out <= 24'h304030;
             12'h344:  out <= 24'h304040;
             12'h345:  out <= 24'h304050;
             12'h346:  out <= 24'h304060;
             12'h347:  out <= 24'h304070;
             12'h348:  out <= 24'h304080;
             12'h349:  out <= 24'h304090;
             12'h34a:  out <= 24'h3040a0;
             12'h34b:  out <= 24'h3040b0;
             12'h34c:  out <= 24'h3040c0;
             12'h34d:  out <= 24'h3040d0;
             12'h34e:  out <= 24'h3040e0;
             12'h34f:  out <= 24'h3040f0;
             12'h350:  out <= 24'h305000;
             12'h351:  out <= 24'h305010;
             12'h352:  out <= 24'h305020;
             12'h353:  out <= 24'h305030;
             12'h354:  out <= 24'h305040;
             12'h355:  out <= 24'h305050;
             12'h356:  out <= 24'h305060;
             12'h357:  out <= 24'h305070;
             12'h358:  out <= 24'h305080;
             12'h359:  out <= 24'h305090;
             12'h35a:  out <= 24'h3050a0;
             12'h35b:  out <= 24'h3050b0;
             12'h35c:  out <= 24'h3050c0;
             12'h35d:  out <= 24'h3050d0;
             12'h35e:  out <= 24'h3050e0;
             12'h35f:  out <= 24'h3050f0;
             12'h360:  out <= 24'h306000;
             12'h361:  out <= 24'h306010;
             12'h362:  out <= 24'h306020;
             12'h363:  out <= 24'h306030;
             12'h364:  out <= 24'h306040;
             12'h365:  out <= 24'h306050;
             12'h366:  out <= 24'h306060;
             12'h367:  out <= 24'h306070;
             12'h368:  out <= 24'h306080;
             12'h369:  out <= 24'h306090;
             12'h36a:  out <= 24'h3060a0;
             12'h36b:  out <= 24'h3060b0;
             12'h36c:  out <= 24'h3060c0;
             12'h36d:  out <= 24'h3060d0;
             12'h36e:  out <= 24'h3060e0;
             12'h36f:  out <= 24'h3060f0;
             12'h370:  out <= 24'h307000;
             12'h371:  out <= 24'h307010;
             12'h372:  out <= 24'h307020;
             12'h373:  out <= 24'h307030;
             12'h374:  out <= 24'h307040;
             12'h375:  out <= 24'h307050;
             12'h376:  out <= 24'h307060;
             12'h377:  out <= 24'h307070;
             12'h378:  out <= 24'h307080;
             12'h379:  out <= 24'h307090;
             12'h37a:  out <= 24'h3070a0;
             12'h37b:  out <= 24'h3070b0;
             12'h37c:  out <= 24'h3070c0;
             12'h37d:  out <= 24'h3070d0;
             12'h37e:  out <= 24'h3070e0;
             12'h37f:  out <= 24'h3070f0;
             12'h380:  out <= 24'h308000;
             12'h381:  out <= 24'h308010;
             12'h382:  out <= 24'h308020;
             12'h383:  out <= 24'h308030;
             12'h384:  out <= 24'h308040;
             12'h385:  out <= 24'h308050;
             12'h386:  out <= 24'h308060;
             12'h387:  out <= 24'h308070;
             12'h388:  out <= 24'h308080;
             12'h389:  out <= 24'h308090;
             12'h38a:  out <= 24'h3080a0;
             12'h38b:  out <= 24'h3080b0;
             12'h38c:  out <= 24'h3080c0;
             12'h38d:  out <= 24'h3080d0;
             12'h38e:  out <= 24'h3080e0;
             12'h38f:  out <= 24'h3080f0;
             12'h390:  out <= 24'h309000;
             12'h391:  out <= 24'h309010;
             12'h392:  out <= 24'h309020;
             12'h393:  out <= 24'h309030;
             12'h394:  out <= 24'h309040;
             12'h395:  out <= 24'h309050;
             12'h396:  out <= 24'h309060;
             12'h397:  out <= 24'h309070;
             12'h398:  out <= 24'h309080;
             12'h399:  out <= 24'h309090;
             12'h39a:  out <= 24'h3090a0;
             12'h39b:  out <= 24'h3090b0;
             12'h39c:  out <= 24'h3090c0;
             12'h39d:  out <= 24'h3090d0;
             12'h39e:  out <= 24'h3090e0;
             12'h39f:  out <= 24'h3090f0;
             12'h3a0:  out <= 24'h30a000;
             12'h3a1:  out <= 24'h30a010;
             12'h3a2:  out <= 24'h30a020;
             12'h3a3:  out <= 24'h30a030;
             12'h3a4:  out <= 24'h30a040;
             12'h3a5:  out <= 24'h30a050;
             12'h3a6:  out <= 24'h30a060;
             12'h3a7:  out <= 24'h30a070;
             12'h3a8:  out <= 24'h30a080;
             12'h3a9:  out <= 24'h30a090;
             12'h3aa:  out <= 24'h30a0a0;
             12'h3ab:  out <= 24'h30a0b0;
             12'h3ac:  out <= 24'h30a0c0;
             12'h3ad:  out <= 24'h30a0d0;
             12'h3ae:  out <= 24'h30a0e0;
             12'h3af:  out <= 24'h30a0f0;
             12'h3b0:  out <= 24'h30b000;
             12'h3b1:  out <= 24'h30b010;
             12'h3b2:  out <= 24'h30b020;
             12'h3b3:  out <= 24'h30b030;
             12'h3b4:  out <= 24'h30b040;
             12'h3b5:  out <= 24'h30b050;
             12'h3b6:  out <= 24'h30b060;
             12'h3b7:  out <= 24'h30b070;
             12'h3b8:  out <= 24'h30b080;
             12'h3b9:  out <= 24'h30b090;
             12'h3ba:  out <= 24'h30b0a0;
             12'h3bb:  out <= 24'h30b0b0;
             12'h3bc:  out <= 24'h30b0c0;
             12'h3bd:  out <= 24'h30b0d0;
             12'h3be:  out <= 24'h30b0e0;
             12'h3bf:  out <= 24'h30b0f0;
             12'h3c0:  out <= 24'h30c000;
             12'h3c1:  out <= 24'h30c010;
             12'h3c2:  out <= 24'h30c020;
             12'h3c3:  out <= 24'h30c030;
             12'h3c4:  out <= 24'h30c040;
             12'h3c5:  out <= 24'h30c050;
             12'h3c6:  out <= 24'h30c060;
             12'h3c7:  out <= 24'h30c070;
             12'h3c8:  out <= 24'h30c080;
             12'h3c9:  out <= 24'h30c090;
             12'h3ca:  out <= 24'h30c0a0;
             12'h3cb:  out <= 24'h30c0b0;
             12'h3cc:  out <= 24'h30c0c0;
             12'h3cd:  out <= 24'h30c0d0;
             12'h3ce:  out <= 24'h30c0e0;
             12'h3cf:  out <= 24'h30c0f0;
             12'h3d0:  out <= 24'h30d000;
             12'h3d1:  out <= 24'h30d010;
             12'h3d2:  out <= 24'h30d020;
             12'h3d3:  out <= 24'h30d030;
             12'h3d4:  out <= 24'h30d040;
             12'h3d5:  out <= 24'h30d050;
             12'h3d6:  out <= 24'h30d060;
             12'h3d7:  out <= 24'h30d070;
             12'h3d8:  out <= 24'h30d080;
             12'h3d9:  out <= 24'h30d090;
             12'h3da:  out <= 24'h30d0a0;
             12'h3db:  out <= 24'h30d0b0;
             12'h3dc:  out <= 24'h30d0c0;
             12'h3dd:  out <= 24'h30d0d0;
             12'h3de:  out <= 24'h30d0e0;
             12'h3df:  out <= 24'h30d0f0;
             12'h3e0:  out <= 24'h30e000;
             12'h3e1:  out <= 24'h30e010;
             12'h3e2:  out <= 24'h30e020;
             12'h3e3:  out <= 24'h30e030;
             12'h3e4:  out <= 24'h30e040;
             12'h3e5:  out <= 24'h30e050;
             12'h3e6:  out <= 24'h30e060;
             12'h3e7:  out <= 24'h30e070;
             12'h3e8:  out <= 24'h30e080;
             12'h3e9:  out <= 24'h30e090;
             12'h3ea:  out <= 24'h30e0a0;
             12'h3eb:  out <= 24'h30e0b0;
             12'h3ec:  out <= 24'h30e0c0;
             12'h3ed:  out <= 24'h30e0d0;
             12'h3ee:  out <= 24'h30e0e0;
             12'h3ef:  out <= 24'h30e0f0;
             12'h3f0:  out <= 24'h30f000;
             12'h3f1:  out <= 24'h30f010;
             12'h3f2:  out <= 24'h30f020;
             12'h3f3:  out <= 24'h30f030;
             12'h3f4:  out <= 24'h30f040;
             12'h3f5:  out <= 24'h30f050;
             12'h3f6:  out <= 24'h30f060;
             12'h3f7:  out <= 24'h30f070;
             12'h3f8:  out <= 24'h30f080;
             12'h3f9:  out <= 24'h30f090;
             12'h3fa:  out <= 24'h30f0a0;
             12'h3fb:  out <= 24'h30f0b0;
             12'h3fc:  out <= 24'h30f0c0;
             12'h3fd:  out <= 24'h30f0d0;
             12'h3fe:  out <= 24'h30f0e0;
             12'h3ff:  out <= 24'h30f0f0;
             12'h400:  out <= 24'h400000;
             12'h401:  out <= 24'h400010;
             12'h402:  out <= 24'h400020;
             12'h403:  out <= 24'h400030;
             12'h404:  out <= 24'h400040;
             12'h405:  out <= 24'h400050;
             12'h406:  out <= 24'h400060;
             12'h407:  out <= 24'h400070;
             12'h408:  out <= 24'h400080;
             12'h409:  out <= 24'h400090;
             12'h40a:  out <= 24'h4000a0;
             12'h40b:  out <= 24'h4000b0;
             12'h40c:  out <= 24'h4000c0;
             12'h40d:  out <= 24'h4000d0;
             12'h40e:  out <= 24'h4000e0;
             12'h40f:  out <= 24'h4000f0;
             12'h410:  out <= 24'h401000;
             12'h411:  out <= 24'h401010;
             12'h412:  out <= 24'h401020;
             12'h413:  out <= 24'h401030;
             12'h414:  out <= 24'h401040;
             12'h415:  out <= 24'h401050;
             12'h416:  out <= 24'h401060;
             12'h417:  out <= 24'h401070;
             12'h418:  out <= 24'h401080;
             12'h419:  out <= 24'h401090;
             12'h41a:  out <= 24'h4010a0;
             12'h41b:  out <= 24'h4010b0;
             12'h41c:  out <= 24'h4010c0;
             12'h41d:  out <= 24'h4010d0;
             12'h41e:  out <= 24'h4010e0;
             12'h41f:  out <= 24'h4010f0;
             12'h420:  out <= 24'h402000;
             12'h421:  out <= 24'h402010;
             12'h422:  out <= 24'h402020;
             12'h423:  out <= 24'h402030;
             12'h424:  out <= 24'h402040;
             12'h425:  out <= 24'h402050;
             12'h426:  out <= 24'h402060;
             12'h427:  out <= 24'h402070;
             12'h428:  out <= 24'h402080;
             12'h429:  out <= 24'h402090;
             12'h42a:  out <= 24'h4020a0;
             12'h42b:  out <= 24'h4020b0;
             12'h42c:  out <= 24'h4020c0;
             12'h42d:  out <= 24'h4020d0;
             12'h42e:  out <= 24'h4020e0;
             12'h42f:  out <= 24'h4020f0;
             12'h430:  out <= 24'h403000;
             12'h431:  out <= 24'h403010;
             12'h432:  out <= 24'h403020;
             12'h433:  out <= 24'h403030;
             12'h434:  out <= 24'h403040;
             12'h435:  out <= 24'h403050;
             12'h436:  out <= 24'h403060;
             12'h437:  out <= 24'h403070;
             12'h438:  out <= 24'h403080;
             12'h439:  out <= 24'h403090;
             12'h43a:  out <= 24'h4030a0;
             12'h43b:  out <= 24'h4030b0;
             12'h43c:  out <= 24'h4030c0;
             12'h43d:  out <= 24'h4030d0;
             12'h43e:  out <= 24'h4030e0;
             12'h43f:  out <= 24'h4030f0;
             12'h440:  out <= 24'h404000;
             12'h441:  out <= 24'h404010;
             12'h442:  out <= 24'h404020;
             12'h443:  out <= 24'h404030;
             12'h444:  out <= 24'h404040;
             12'h445:  out <= 24'h404050;
             12'h446:  out <= 24'h404060;
             12'h447:  out <= 24'h404070;
             12'h448:  out <= 24'h404080;
             12'h449:  out <= 24'h404090;
             12'h44a:  out <= 24'h4040a0;
             12'h44b:  out <= 24'h4040b0;
             12'h44c:  out <= 24'h4040c0;
             12'h44d:  out <= 24'h4040d0;
             12'h44e:  out <= 24'h4040e0;
             12'h44f:  out <= 24'h4040f0;
             12'h450:  out <= 24'h405000;
             12'h451:  out <= 24'h405010;
             12'h452:  out <= 24'h405020;
             12'h453:  out <= 24'h405030;
             12'h454:  out <= 24'h405040;
             12'h455:  out <= 24'h405050;
             12'h456:  out <= 24'h405060;
             12'h457:  out <= 24'h405070;
             12'h458:  out <= 24'h405080;
             12'h459:  out <= 24'h405090;
             12'h45a:  out <= 24'h4050a0;
             12'h45b:  out <= 24'h4050b0;
             12'h45c:  out <= 24'h4050c0;
             12'h45d:  out <= 24'h4050d0;
             12'h45e:  out <= 24'h4050e0;
             12'h45f:  out <= 24'h4050f0;
             12'h460:  out <= 24'h406000;
             12'h461:  out <= 24'h406010;
             12'h462:  out <= 24'h406020;
             12'h463:  out <= 24'h406030;
             12'h464:  out <= 24'h406040;
             12'h465:  out <= 24'h406050;
             12'h466:  out <= 24'h406060;
             12'h467:  out <= 24'h406070;
             12'h468:  out <= 24'h406080;
             12'h469:  out <= 24'h406090;
             12'h46a:  out <= 24'h4060a0;
             12'h46b:  out <= 24'h4060b0;
             12'h46c:  out <= 24'h4060c0;
             12'h46d:  out <= 24'h4060d0;
             12'h46e:  out <= 24'h4060e0;
             12'h46f:  out <= 24'h4060f0;
             12'h470:  out <= 24'h407000;
             12'h471:  out <= 24'h407010;
             12'h472:  out <= 24'h407020;
             12'h473:  out <= 24'h407030;
             12'h474:  out <= 24'h407040;
             12'h475:  out <= 24'h407050;
             12'h476:  out <= 24'h407060;
             12'h477:  out <= 24'h407070;
             12'h478:  out <= 24'h407080;
             12'h479:  out <= 24'h407090;
             12'h47a:  out <= 24'h4070a0;
             12'h47b:  out <= 24'h4070b0;
             12'h47c:  out <= 24'h4070c0;
             12'h47d:  out <= 24'h4070d0;
             12'h47e:  out <= 24'h4070e0;
             12'h47f:  out <= 24'h4070f0;
             12'h480:  out <= 24'h408000;
             12'h481:  out <= 24'h408010;
             12'h482:  out <= 24'h408020;
             12'h483:  out <= 24'h408030;
             12'h484:  out <= 24'h408040;
             12'h485:  out <= 24'h408050;
             12'h486:  out <= 24'h408060;
             12'h487:  out <= 24'h408070;
             12'h488:  out <= 24'h408080;
             12'h489:  out <= 24'h408090;
             12'h48a:  out <= 24'h4080a0;
             12'h48b:  out <= 24'h4080b0;
             12'h48c:  out <= 24'h4080c0;
             12'h48d:  out <= 24'h4080d0;
             12'h48e:  out <= 24'h4080e0;
             12'h48f:  out <= 24'h4080f0;
             12'h490:  out <= 24'h409000;
             12'h491:  out <= 24'h409010;
             12'h492:  out <= 24'h409020;
             12'h493:  out <= 24'h409030;
             12'h494:  out <= 24'h409040;
             12'h495:  out <= 24'h409050;
             12'h496:  out <= 24'h409060;
             12'h497:  out <= 24'h409070;
             12'h498:  out <= 24'h409080;
             12'h499:  out <= 24'h409090;
             12'h49a:  out <= 24'h4090a0;
             12'h49b:  out <= 24'h4090b0;
             12'h49c:  out <= 24'h4090c0;
             12'h49d:  out <= 24'h4090d0;
             12'h49e:  out <= 24'h4090e0;
             12'h49f:  out <= 24'h4090f0;
             12'h4a0:  out <= 24'h40a000;
             12'h4a1:  out <= 24'h40a010;
             12'h4a2:  out <= 24'h40a020;
             12'h4a3:  out <= 24'h40a030;
             12'h4a4:  out <= 24'h40a040;
             12'h4a5:  out <= 24'h40a050;
             12'h4a6:  out <= 24'h40a060;
             12'h4a7:  out <= 24'h40a070;
             12'h4a8:  out <= 24'h40a080;
             12'h4a9:  out <= 24'h40a090;
             12'h4aa:  out <= 24'h40a0a0;
             12'h4ab:  out <= 24'h40a0b0;
             12'h4ac:  out <= 24'h40a0c0;
             12'h4ad:  out <= 24'h40a0d0;
             12'h4ae:  out <= 24'h40a0e0;
             12'h4af:  out <= 24'h40a0f0;
             12'h4b0:  out <= 24'h40b000;
             12'h4b1:  out <= 24'h40b010;
             12'h4b2:  out <= 24'h40b020;
             12'h4b3:  out <= 24'h40b030;
             12'h4b4:  out <= 24'h40b040;
             12'h4b5:  out <= 24'h40b050;
             12'h4b6:  out <= 24'h40b060;
             12'h4b7:  out <= 24'h40b070;
             12'h4b8:  out <= 24'h40b080;
             12'h4b9:  out <= 24'h40b090;
             12'h4ba:  out <= 24'h40b0a0;
             12'h4bb:  out <= 24'h40b0b0;
             12'h4bc:  out <= 24'h40b0c0;
             12'h4bd:  out <= 24'h40b0d0;
             12'h4be:  out <= 24'h40b0e0;
             12'h4bf:  out <= 24'h40b0f0;
             12'h4c0:  out <= 24'h40c000;
             12'h4c1:  out <= 24'h40c010;
             12'h4c2:  out <= 24'h40c020;
             12'h4c3:  out <= 24'h40c030;
             12'h4c4:  out <= 24'h40c040;
             12'h4c5:  out <= 24'h40c050;
             12'h4c6:  out <= 24'h40c060;
             12'h4c7:  out <= 24'h40c070;
             12'h4c8:  out <= 24'h40c080;
             12'h4c9:  out <= 24'h40c090;
             12'h4ca:  out <= 24'h40c0a0;
             12'h4cb:  out <= 24'h40c0b0;
             12'h4cc:  out <= 24'h40c0c0;
             12'h4cd:  out <= 24'h40c0d0;
             12'h4ce:  out <= 24'h40c0e0;
             12'h4cf:  out <= 24'h40c0f0;
             12'h4d0:  out <= 24'h40d000;
             12'h4d1:  out <= 24'h40d010;
             12'h4d2:  out <= 24'h40d020;
             12'h4d3:  out <= 24'h40d030;
             12'h4d4:  out <= 24'h40d040;
             12'h4d5:  out <= 24'h40d050;
             12'h4d6:  out <= 24'h40d060;
             12'h4d7:  out <= 24'h40d070;
             12'h4d8:  out <= 24'h40d080;
             12'h4d9:  out <= 24'h40d090;
             12'h4da:  out <= 24'h40d0a0;
             12'h4db:  out <= 24'h40d0b0;
             12'h4dc:  out <= 24'h40d0c0;
             12'h4dd:  out <= 24'h40d0d0;
             12'h4de:  out <= 24'h40d0e0;
             12'h4df:  out <= 24'h40d0f0;
             12'h4e0:  out <= 24'h40e000;
             12'h4e1:  out <= 24'h40e010;
             12'h4e2:  out <= 24'h40e020;
             12'h4e3:  out <= 24'h40e030;
             12'h4e4:  out <= 24'h40e040;
             12'h4e5:  out <= 24'h40e050;
             12'h4e6:  out <= 24'h40e060;
             12'h4e7:  out <= 24'h40e070;
             12'h4e8:  out <= 24'h40e080;
             12'h4e9:  out <= 24'h40e090;
             12'h4ea:  out <= 24'h40e0a0;
             12'h4eb:  out <= 24'h40e0b0;
             12'h4ec:  out <= 24'h40e0c0;
             12'h4ed:  out <= 24'h40e0d0;
             12'h4ee:  out <= 24'h40e0e0;
             12'h4ef:  out <= 24'h40e0f0;
             12'h4f0:  out <= 24'h40f000;
             12'h4f1:  out <= 24'h40f010;
             12'h4f2:  out <= 24'h40f020;
             12'h4f3:  out <= 24'h40f030;
             12'h4f4:  out <= 24'h40f040;
             12'h4f5:  out <= 24'h40f050;
             12'h4f6:  out <= 24'h40f060;
             12'h4f7:  out <= 24'h40f070;
             12'h4f8:  out <= 24'h40f080;
             12'h4f9:  out <= 24'h40f090;
             12'h4fa:  out <= 24'h40f0a0;
             12'h4fb:  out <= 24'h40f0b0;
             12'h4fc:  out <= 24'h40f0c0;
             12'h4fd:  out <= 24'h40f0d0;
             12'h4fe:  out <= 24'h40f0e0;
             12'h4ff:  out <= 24'h40f0f0;
             12'h500:  out <= 24'h500000;
             12'h501:  out <= 24'h500010;
             12'h502:  out <= 24'h500020;
             12'h503:  out <= 24'h500030;
             12'h504:  out <= 24'h500040;
             12'h505:  out <= 24'h500050;
             12'h506:  out <= 24'h500060;
             12'h507:  out <= 24'h500070;
             12'h508:  out <= 24'h500080;
             12'h509:  out <= 24'h500090;
             12'h50a:  out <= 24'h5000a0;
             12'h50b:  out <= 24'h5000b0;
             12'h50c:  out <= 24'h5000c0;
             12'h50d:  out <= 24'h5000d0;
             12'h50e:  out <= 24'h5000e0;
             12'h50f:  out <= 24'h5000f0;
             12'h510:  out <= 24'h501000;
             12'h511:  out <= 24'h501010;
             12'h512:  out <= 24'h501020;
             12'h513:  out <= 24'h501030;
             12'h514:  out <= 24'h501040;
             12'h515:  out <= 24'h501050;
             12'h516:  out <= 24'h501060;
             12'h517:  out <= 24'h501070;
             12'h518:  out <= 24'h501080;
             12'h519:  out <= 24'h501090;
             12'h51a:  out <= 24'h5010a0;
             12'h51b:  out <= 24'h5010b0;
             12'h51c:  out <= 24'h5010c0;
             12'h51d:  out <= 24'h5010d0;
             12'h51e:  out <= 24'h5010e0;
             12'h51f:  out <= 24'h5010f0;
             12'h520:  out <= 24'h502000;
             12'h521:  out <= 24'h502010;
             12'h522:  out <= 24'h502020;
             12'h523:  out <= 24'h502030;
             12'h524:  out <= 24'h502040;
             12'h525:  out <= 24'h502050;
             12'h526:  out <= 24'h502060;
             12'h527:  out <= 24'h502070;
             12'h528:  out <= 24'h502080;
             12'h529:  out <= 24'h502090;
             12'h52a:  out <= 24'h5020a0;
             12'h52b:  out <= 24'h5020b0;
             12'h52c:  out <= 24'h5020c0;
             12'h52d:  out <= 24'h5020d0;
             12'h52e:  out <= 24'h5020e0;
             12'h52f:  out <= 24'h5020f0;
             12'h530:  out <= 24'h503000;
             12'h531:  out <= 24'h503010;
             12'h532:  out <= 24'h503020;
             12'h533:  out <= 24'h503030;
             12'h534:  out <= 24'h503040;
             12'h535:  out <= 24'h503050;
             12'h536:  out <= 24'h503060;
             12'h537:  out <= 24'h503070;
             12'h538:  out <= 24'h503080;
             12'h539:  out <= 24'h503090;
             12'h53a:  out <= 24'h5030a0;
             12'h53b:  out <= 24'h5030b0;
             12'h53c:  out <= 24'h5030c0;
             12'h53d:  out <= 24'h5030d0;
             12'h53e:  out <= 24'h5030e0;
             12'h53f:  out <= 24'h5030f0;
             12'h540:  out <= 24'h504000;
             12'h541:  out <= 24'h504010;
             12'h542:  out <= 24'h504020;
             12'h543:  out <= 24'h504030;
             12'h544:  out <= 24'h504040;
             12'h545:  out <= 24'h504050;
             12'h546:  out <= 24'h504060;
             12'h547:  out <= 24'h504070;
             12'h548:  out <= 24'h504080;
             12'h549:  out <= 24'h504090;
             12'h54a:  out <= 24'h5040a0;
             12'h54b:  out <= 24'h5040b0;
             12'h54c:  out <= 24'h5040c0;
             12'h54d:  out <= 24'h5040d0;
             12'h54e:  out <= 24'h5040e0;
             12'h54f:  out <= 24'h5040f0;
             12'h550:  out <= 24'h505000;
             12'h551:  out <= 24'h505010;
             12'h552:  out <= 24'h505020;
             12'h553:  out <= 24'h505030;
             12'h554:  out <= 24'h505040;
             12'h555:  out <= 24'h505050;
             12'h556:  out <= 24'h505060;
             12'h557:  out <= 24'h505070;
             12'h558:  out <= 24'h505080;
             12'h559:  out <= 24'h505090;
             12'h55a:  out <= 24'h5050a0;
             12'h55b:  out <= 24'h5050b0;
             12'h55c:  out <= 24'h5050c0;
             12'h55d:  out <= 24'h5050d0;
             12'h55e:  out <= 24'h5050e0;
             12'h55f:  out <= 24'h5050f0;
             12'h560:  out <= 24'h506000;
             12'h561:  out <= 24'h506010;
             12'h562:  out <= 24'h506020;
             12'h563:  out <= 24'h506030;
             12'h564:  out <= 24'h506040;
             12'h565:  out <= 24'h506050;
             12'h566:  out <= 24'h506060;
             12'h567:  out <= 24'h506070;
             12'h568:  out <= 24'h506080;
             12'h569:  out <= 24'h506090;
             12'h56a:  out <= 24'h5060a0;
             12'h56b:  out <= 24'h5060b0;
             12'h56c:  out <= 24'h5060c0;
             12'h56d:  out <= 24'h5060d0;
             12'h56e:  out <= 24'h5060e0;
             12'h56f:  out <= 24'h5060f0;
             12'h570:  out <= 24'h507000;
             12'h571:  out <= 24'h507010;
             12'h572:  out <= 24'h507020;
             12'h573:  out <= 24'h507030;
             12'h574:  out <= 24'h507040;
             12'h575:  out <= 24'h507050;
             12'h576:  out <= 24'h507060;
             12'h577:  out <= 24'h507070;
             12'h578:  out <= 24'h507080;
             12'h579:  out <= 24'h507090;
             12'h57a:  out <= 24'h5070a0;
             12'h57b:  out <= 24'h5070b0;
             12'h57c:  out <= 24'h5070c0;
             12'h57d:  out <= 24'h5070d0;
             12'h57e:  out <= 24'h5070e0;
             12'h57f:  out <= 24'h5070f0;
             12'h580:  out <= 24'h508000;
             12'h581:  out <= 24'h508010;
             12'h582:  out <= 24'h508020;
             12'h583:  out <= 24'h508030;
             12'h584:  out <= 24'h508040;
             12'h585:  out <= 24'h508050;
             12'h586:  out <= 24'h508060;
             12'h587:  out <= 24'h508070;
             12'h588:  out <= 24'h508080;
             12'h589:  out <= 24'h508090;
             12'h58a:  out <= 24'h5080a0;
             12'h58b:  out <= 24'h5080b0;
             12'h58c:  out <= 24'h5080c0;
             12'h58d:  out <= 24'h5080d0;
             12'h58e:  out <= 24'h5080e0;
             12'h58f:  out <= 24'h5080f0;
             12'h590:  out <= 24'h509000;
             12'h591:  out <= 24'h509010;
             12'h592:  out <= 24'h509020;
             12'h593:  out <= 24'h509030;
             12'h594:  out <= 24'h509040;
             12'h595:  out <= 24'h509050;
             12'h596:  out <= 24'h509060;
             12'h597:  out <= 24'h509070;
             12'h598:  out <= 24'h509080;
             12'h599:  out <= 24'h509090;
             12'h59a:  out <= 24'h5090a0;
             12'h59b:  out <= 24'h5090b0;
             12'h59c:  out <= 24'h5090c0;
             12'h59d:  out <= 24'h5090d0;
             12'h59e:  out <= 24'h5090e0;
             12'h59f:  out <= 24'h5090f0;
             12'h5a0:  out <= 24'h50a000;
             12'h5a1:  out <= 24'h50a010;
             12'h5a2:  out <= 24'h50a020;
             12'h5a3:  out <= 24'h50a030;
             12'h5a4:  out <= 24'h50a040;
             12'h5a5:  out <= 24'h50a050;
             12'h5a6:  out <= 24'h50a060;
             12'h5a7:  out <= 24'h50a070;
             12'h5a8:  out <= 24'h50a080;
             12'h5a9:  out <= 24'h50a090;
             12'h5aa:  out <= 24'h50a0a0;
             12'h5ab:  out <= 24'h50a0b0;
             12'h5ac:  out <= 24'h50a0c0;
             12'h5ad:  out <= 24'h50a0d0;
             12'h5ae:  out <= 24'h50a0e0;
             12'h5af:  out <= 24'h50a0f0;
             12'h5b0:  out <= 24'h50b000;
             12'h5b1:  out <= 24'h50b010;
             12'h5b2:  out <= 24'h50b020;
             12'h5b3:  out <= 24'h50b030;
             12'h5b4:  out <= 24'h50b040;
             12'h5b5:  out <= 24'h50b050;
             12'h5b6:  out <= 24'h50b060;
             12'h5b7:  out <= 24'h50b070;
             12'h5b8:  out <= 24'h50b080;
             12'h5b9:  out <= 24'h50b090;
             12'h5ba:  out <= 24'h50b0a0;
             12'h5bb:  out <= 24'h50b0b0;
             12'h5bc:  out <= 24'h50b0c0;
             12'h5bd:  out <= 24'h50b0d0;
             12'h5be:  out <= 24'h50b0e0;
             12'h5bf:  out <= 24'h50b0f0;
             12'h5c0:  out <= 24'h50c000;
             12'h5c1:  out <= 24'h50c010;
             12'h5c2:  out <= 24'h50c020;
             12'h5c3:  out <= 24'h50c030;
             12'h5c4:  out <= 24'h50c040;
             12'h5c5:  out <= 24'h50c050;
             12'h5c6:  out <= 24'h50c060;
             12'h5c7:  out <= 24'h50c070;
             12'h5c8:  out <= 24'h50c080;
             12'h5c9:  out <= 24'h50c090;
             12'h5ca:  out <= 24'h50c0a0;
             12'h5cb:  out <= 24'h50c0b0;
             12'h5cc:  out <= 24'h50c0c0;
             12'h5cd:  out <= 24'h50c0d0;
             12'h5ce:  out <= 24'h50c0e0;
             12'h5cf:  out <= 24'h50c0f0;
             12'h5d0:  out <= 24'h50d000;
             12'h5d1:  out <= 24'h50d010;
             12'h5d2:  out <= 24'h50d020;
             12'h5d3:  out <= 24'h50d030;
             12'h5d4:  out <= 24'h50d040;
             12'h5d5:  out <= 24'h50d050;
             12'h5d6:  out <= 24'h50d060;
             12'h5d7:  out <= 24'h50d070;
             12'h5d8:  out <= 24'h50d080;
             12'h5d9:  out <= 24'h50d090;
             12'h5da:  out <= 24'h50d0a0;
             12'h5db:  out <= 24'h50d0b0;
             12'h5dc:  out <= 24'h50d0c0;
             12'h5dd:  out <= 24'h50d0d0;
             12'h5de:  out <= 24'h50d0e0;
             12'h5df:  out <= 24'h50d0f0;
             12'h5e0:  out <= 24'h50e000;
             12'h5e1:  out <= 24'h50e010;
             12'h5e2:  out <= 24'h50e020;
             12'h5e3:  out <= 24'h50e030;
             12'h5e4:  out <= 24'h50e040;
             12'h5e5:  out <= 24'h50e050;
             12'h5e6:  out <= 24'h50e060;
             12'h5e7:  out <= 24'h50e070;
             12'h5e8:  out <= 24'h50e080;
             12'h5e9:  out <= 24'h50e090;
             12'h5ea:  out <= 24'h50e0a0;
             12'h5eb:  out <= 24'h50e0b0;
             12'h5ec:  out <= 24'h50e0c0;
             12'h5ed:  out <= 24'h50e0d0;
             12'h5ee:  out <= 24'h50e0e0;
             12'h5ef:  out <= 24'h50e0f0;
             12'h5f0:  out <= 24'h50f000;
             12'h5f1:  out <= 24'h50f010;
             12'h5f2:  out <= 24'h50f020;
             12'h5f3:  out <= 24'h50f030;
             12'h5f4:  out <= 24'h50f040;
             12'h5f5:  out <= 24'h50f050;
             12'h5f6:  out <= 24'h50f060;
             12'h5f7:  out <= 24'h50f070;
             12'h5f8:  out <= 24'h50f080;
             12'h5f9:  out <= 24'h50f090;
             12'h5fa:  out <= 24'h50f0a0;
             12'h5fb:  out <= 24'h50f0b0;
             12'h5fc:  out <= 24'h50f0c0;
             12'h5fd:  out <= 24'h50f0d0;
             12'h5fe:  out <= 24'h50f0e0;
             12'h5ff:  out <= 24'h50f0f0;
             12'h600:  out <= 24'h600000;
             12'h601:  out <= 24'h600010;
             12'h602:  out <= 24'h600020;
             12'h603:  out <= 24'h600030;
             12'h604:  out <= 24'h600040;
             12'h605:  out <= 24'h600050;
             12'h606:  out <= 24'h600060;
             12'h607:  out <= 24'h600070;
             12'h608:  out <= 24'h600080;
             12'h609:  out <= 24'h600090;
             12'h60a:  out <= 24'h6000a0;
             12'h60b:  out <= 24'h6000b0;
             12'h60c:  out <= 24'h6000c0;
             12'h60d:  out <= 24'h6000d0;
             12'h60e:  out <= 24'h6000e0;
             12'h60f:  out <= 24'h6000f0;
             12'h610:  out <= 24'h601000;
             12'h611:  out <= 24'h601010;
             12'h612:  out <= 24'h601020;
             12'h613:  out <= 24'h601030;
             12'h614:  out <= 24'h601040;
             12'h615:  out <= 24'h601050;
             12'h616:  out <= 24'h601060;
             12'h617:  out <= 24'h601070;
             12'h618:  out <= 24'h601080;
             12'h619:  out <= 24'h601090;
             12'h61a:  out <= 24'h6010a0;
             12'h61b:  out <= 24'h6010b0;
             12'h61c:  out <= 24'h6010c0;
             12'h61d:  out <= 24'h6010d0;
             12'h61e:  out <= 24'h6010e0;
             12'h61f:  out <= 24'h6010f0;
             12'h620:  out <= 24'h602000;
             12'h621:  out <= 24'h602010;
             12'h622:  out <= 24'h602020;
             12'h623:  out <= 24'h602030;
             12'h624:  out <= 24'h602040;
             12'h625:  out <= 24'h602050;
             12'h626:  out <= 24'h602060;
             12'h627:  out <= 24'h602070;
             12'h628:  out <= 24'h602080;
             12'h629:  out <= 24'h602090;
             12'h62a:  out <= 24'h6020a0;
             12'h62b:  out <= 24'h6020b0;
             12'h62c:  out <= 24'h6020c0;
             12'h62d:  out <= 24'h6020d0;
             12'h62e:  out <= 24'h6020e0;
             12'h62f:  out <= 24'h6020f0;
             12'h630:  out <= 24'h603000;
             12'h631:  out <= 24'h603010;
             12'h632:  out <= 24'h603020;
             12'h633:  out <= 24'h603030;
             12'h634:  out <= 24'h603040;
             12'h635:  out <= 24'h603050;
             12'h636:  out <= 24'h603060;
             12'h637:  out <= 24'h603070;
             12'h638:  out <= 24'h603080;
             12'h639:  out <= 24'h603090;
             12'h63a:  out <= 24'h6030a0;
             12'h63b:  out <= 24'h6030b0;
             12'h63c:  out <= 24'h6030c0;
             12'h63d:  out <= 24'h6030d0;
             12'h63e:  out <= 24'h6030e0;
             12'h63f:  out <= 24'h6030f0;
             12'h640:  out <= 24'h604000;
             12'h641:  out <= 24'h604010;
             12'h642:  out <= 24'h604020;
             12'h643:  out <= 24'h604030;
             12'h644:  out <= 24'h604040;
             12'h645:  out <= 24'h604050;
             12'h646:  out <= 24'h604060;
             12'h647:  out <= 24'h604070;
             12'h648:  out <= 24'h604080;
             12'h649:  out <= 24'h604090;
             12'h64a:  out <= 24'h6040a0;
             12'h64b:  out <= 24'h6040b0;
             12'h64c:  out <= 24'h6040c0;
             12'h64d:  out <= 24'h6040d0;
             12'h64e:  out <= 24'h6040e0;
             12'h64f:  out <= 24'h6040f0;
             12'h650:  out <= 24'h605000;
             12'h651:  out <= 24'h605010;
             12'h652:  out <= 24'h605020;
             12'h653:  out <= 24'h605030;
             12'h654:  out <= 24'h605040;
             12'h655:  out <= 24'h605050;
             12'h656:  out <= 24'h605060;
             12'h657:  out <= 24'h605070;
             12'h658:  out <= 24'h605080;
             12'h659:  out <= 24'h605090;
             12'h65a:  out <= 24'h6050a0;
             12'h65b:  out <= 24'h6050b0;
             12'h65c:  out <= 24'h6050c0;
             12'h65d:  out <= 24'h6050d0;
             12'h65e:  out <= 24'h6050e0;
             12'h65f:  out <= 24'h6050f0;
             12'h660:  out <= 24'h606000;
             12'h661:  out <= 24'h606010;
             12'h662:  out <= 24'h606020;
             12'h663:  out <= 24'h606030;
             12'h664:  out <= 24'h606040;
             12'h665:  out <= 24'h606050;
             12'h666:  out <= 24'h606060;
             12'h667:  out <= 24'h606070;
             12'h668:  out <= 24'h606080;
             12'h669:  out <= 24'h606090;
             12'h66a:  out <= 24'h6060a0;
             12'h66b:  out <= 24'h6060b0;
             12'h66c:  out <= 24'h6060c0;
             12'h66d:  out <= 24'h6060d0;
             12'h66e:  out <= 24'h6060e0;
             12'h66f:  out <= 24'h6060f0;
             12'h670:  out <= 24'h607000;
             12'h671:  out <= 24'h607010;
             12'h672:  out <= 24'h607020;
             12'h673:  out <= 24'h607030;
             12'h674:  out <= 24'h607040;
             12'h675:  out <= 24'h607050;
             12'h676:  out <= 24'h607060;
             12'h677:  out <= 24'h607070;
             12'h678:  out <= 24'h607080;
             12'h679:  out <= 24'h607090;
             12'h67a:  out <= 24'h6070a0;
             12'h67b:  out <= 24'h6070b0;
             12'h67c:  out <= 24'h6070c0;
             12'h67d:  out <= 24'h6070d0;
             12'h67e:  out <= 24'h6070e0;
             12'h67f:  out <= 24'h6070f0;
             12'h680:  out <= 24'h608000;
             12'h681:  out <= 24'h608010;
             12'h682:  out <= 24'h608020;
             12'h683:  out <= 24'h608030;
             12'h684:  out <= 24'h608040;
             12'h685:  out <= 24'h608050;
             12'h686:  out <= 24'h608060;
             12'h687:  out <= 24'h608070;
             12'h688:  out <= 24'h608080;
             12'h689:  out <= 24'h608090;
             12'h68a:  out <= 24'h6080a0;
             12'h68b:  out <= 24'h6080b0;
             12'h68c:  out <= 24'h6080c0;
             12'h68d:  out <= 24'h6080d0;
             12'h68e:  out <= 24'h6080e0;
             12'h68f:  out <= 24'h6080f0;
             12'h690:  out <= 24'h609000;
             12'h691:  out <= 24'h609010;
             12'h692:  out <= 24'h609020;
             12'h693:  out <= 24'h609030;
             12'h694:  out <= 24'h609040;
             12'h695:  out <= 24'h609050;
             12'h696:  out <= 24'h609060;
             12'h697:  out <= 24'h609070;
             12'h698:  out <= 24'h609080;
             12'h699:  out <= 24'h609090;
             12'h69a:  out <= 24'h6090a0;
             12'h69b:  out <= 24'h6090b0;
             12'h69c:  out <= 24'h6090c0;
             12'h69d:  out <= 24'h6090d0;
             12'h69e:  out <= 24'h6090e0;
             12'h69f:  out <= 24'h6090f0;
             12'h6a0:  out <= 24'h60a000;
             12'h6a1:  out <= 24'h60a010;
             12'h6a2:  out <= 24'h60a020;
             12'h6a3:  out <= 24'h60a030;
             12'h6a4:  out <= 24'h60a040;
             12'h6a5:  out <= 24'h60a050;
             12'h6a6:  out <= 24'h60a060;
             12'h6a7:  out <= 24'h60a070;
             12'h6a8:  out <= 24'h60a080;
             12'h6a9:  out <= 24'h60a090;
             12'h6aa:  out <= 24'h60a0a0;
             12'h6ab:  out <= 24'h60a0b0;
             12'h6ac:  out <= 24'h60a0c0;
             12'h6ad:  out <= 24'h60a0d0;
             12'h6ae:  out <= 24'h60a0e0;
             12'h6af:  out <= 24'h60a0f0;
             12'h6b0:  out <= 24'h60b000;
             12'h6b1:  out <= 24'h60b010;
             12'h6b2:  out <= 24'h60b020;
             12'h6b3:  out <= 24'h60b030;
             12'h6b4:  out <= 24'h60b040;
             12'h6b5:  out <= 24'h60b050;
             12'h6b6:  out <= 24'h60b060;
             12'h6b7:  out <= 24'h60b070;
             12'h6b8:  out <= 24'h60b080;
             12'h6b9:  out <= 24'h60b090;
             12'h6ba:  out <= 24'h60b0a0;
             12'h6bb:  out <= 24'h60b0b0;
             12'h6bc:  out <= 24'h60b0c0;
             12'h6bd:  out <= 24'h60b0d0;
             12'h6be:  out <= 24'h60b0e0;
             12'h6bf:  out <= 24'h60b0f0;
             12'h6c0:  out <= 24'h60c000;
             12'h6c1:  out <= 24'h60c010;
             12'h6c2:  out <= 24'h60c020;
             12'h6c3:  out <= 24'h60c030;
             12'h6c4:  out <= 24'h60c040;
             12'h6c5:  out <= 24'h60c050;
             12'h6c6:  out <= 24'h60c060;
             12'h6c7:  out <= 24'h60c070;
             12'h6c8:  out <= 24'h60c080;
             12'h6c9:  out <= 24'h60c090;
             12'h6ca:  out <= 24'h60c0a0;
             12'h6cb:  out <= 24'h60c0b0;
             12'h6cc:  out <= 24'h60c0c0;
             12'h6cd:  out <= 24'h60c0d0;
             12'h6ce:  out <= 24'h60c0e0;
             12'h6cf:  out <= 24'h60c0f0;
             12'h6d0:  out <= 24'h60d000;
             12'h6d1:  out <= 24'h60d010;
             12'h6d2:  out <= 24'h60d020;
             12'h6d3:  out <= 24'h60d030;
             12'h6d4:  out <= 24'h60d040;
             12'h6d5:  out <= 24'h60d050;
             12'h6d6:  out <= 24'h60d060;
             12'h6d7:  out <= 24'h60d070;
             12'h6d8:  out <= 24'h60d080;
             12'h6d9:  out <= 24'h60d090;
             12'h6da:  out <= 24'h60d0a0;
             12'h6db:  out <= 24'h60d0b0;
             12'h6dc:  out <= 24'h60d0c0;
             12'h6dd:  out <= 24'h60d0d0;
             12'h6de:  out <= 24'h60d0e0;
             12'h6df:  out <= 24'h60d0f0;
             12'h6e0:  out <= 24'h60e000;
             12'h6e1:  out <= 24'h60e010;
             12'h6e2:  out <= 24'h60e020;
             12'h6e3:  out <= 24'h60e030;
             12'h6e4:  out <= 24'h60e040;
             12'h6e5:  out <= 24'h60e050;
             12'h6e6:  out <= 24'h60e060;
             12'h6e7:  out <= 24'h60e070;
             12'h6e8:  out <= 24'h60e080;
             12'h6e9:  out <= 24'h60e090;
             12'h6ea:  out <= 24'h60e0a0;
             12'h6eb:  out <= 24'h60e0b0;
             12'h6ec:  out <= 24'h60e0c0;
             12'h6ed:  out <= 24'h60e0d0;
             12'h6ee:  out <= 24'h60e0e0;
             12'h6ef:  out <= 24'h60e0f0;
             12'h6f0:  out <= 24'h60f000;
             12'h6f1:  out <= 24'h60f010;
             12'h6f2:  out <= 24'h60f020;
             12'h6f3:  out <= 24'h60f030;
             12'h6f4:  out <= 24'h60f040;
             12'h6f5:  out <= 24'h60f050;
             12'h6f6:  out <= 24'h60f060;
             12'h6f7:  out <= 24'h60f070;
             12'h6f8:  out <= 24'h60f080;
             12'h6f9:  out <= 24'h60f090;
             12'h6fa:  out <= 24'h60f0a0;
             12'h6fb:  out <= 24'h60f0b0;
             12'h6fc:  out <= 24'h60f0c0;
             12'h6fd:  out <= 24'h60f0d0;
             12'h6fe:  out <= 24'h60f0e0;
             12'h6ff:  out <= 24'h60f0f0;
             12'h700:  out <= 24'h700000;
             12'h701:  out <= 24'h700010;
             12'h702:  out <= 24'h700020;
             12'h703:  out <= 24'h700030;
             12'h704:  out <= 24'h700040;
             12'h705:  out <= 24'h700050;
             12'h706:  out <= 24'h700060;
             12'h707:  out <= 24'h700070;
             12'h708:  out <= 24'h700080;
             12'h709:  out <= 24'h700090;
             12'h70a:  out <= 24'h7000a0;
             12'h70b:  out <= 24'h7000b0;
             12'h70c:  out <= 24'h7000c0;
             12'h70d:  out <= 24'h7000d0;
             12'h70e:  out <= 24'h7000e0;
             12'h70f:  out <= 24'h7000f0;
             12'h710:  out <= 24'h701000;
             12'h711:  out <= 24'h701010;
             12'h712:  out <= 24'h701020;
             12'h713:  out <= 24'h701030;
             12'h714:  out <= 24'h701040;
             12'h715:  out <= 24'h701050;
             12'h716:  out <= 24'h701060;
             12'h717:  out <= 24'h701070;
             12'h718:  out <= 24'h701080;
             12'h719:  out <= 24'h701090;
             12'h71a:  out <= 24'h7010a0;
             12'h71b:  out <= 24'h7010b0;
             12'h71c:  out <= 24'h7010c0;
             12'h71d:  out <= 24'h7010d0;
             12'h71e:  out <= 24'h7010e0;
             12'h71f:  out <= 24'h7010f0;
             12'h720:  out <= 24'h702000;
             12'h721:  out <= 24'h702010;
             12'h722:  out <= 24'h702020;
             12'h723:  out <= 24'h702030;
             12'h724:  out <= 24'h702040;
             12'h725:  out <= 24'h702050;
             12'h726:  out <= 24'h702060;
             12'h727:  out <= 24'h702070;
             12'h728:  out <= 24'h702080;
             12'h729:  out <= 24'h702090;
             12'h72a:  out <= 24'h7020a0;
             12'h72b:  out <= 24'h7020b0;
             12'h72c:  out <= 24'h7020c0;
             12'h72d:  out <= 24'h7020d0;
             12'h72e:  out <= 24'h7020e0;
             12'h72f:  out <= 24'h7020f0;
             12'h730:  out <= 24'h703000;
             12'h731:  out <= 24'h703010;
             12'h732:  out <= 24'h703020;
             12'h733:  out <= 24'h703030;
             12'h734:  out <= 24'h703040;
             12'h735:  out <= 24'h703050;
             12'h736:  out <= 24'h703060;
             12'h737:  out <= 24'h703070;
             12'h738:  out <= 24'h703080;
             12'h739:  out <= 24'h703090;
             12'h73a:  out <= 24'h7030a0;
             12'h73b:  out <= 24'h7030b0;
             12'h73c:  out <= 24'h7030c0;
             12'h73d:  out <= 24'h7030d0;
             12'h73e:  out <= 24'h7030e0;
             12'h73f:  out <= 24'h7030f0;
             12'h740:  out <= 24'h704000;
             12'h741:  out <= 24'h704010;
             12'h742:  out <= 24'h704020;
             12'h743:  out <= 24'h704030;
             12'h744:  out <= 24'h704040;
             12'h745:  out <= 24'h704050;
             12'h746:  out <= 24'h704060;
             12'h747:  out <= 24'h704070;
             12'h748:  out <= 24'h704080;
             12'h749:  out <= 24'h704090;
             12'h74a:  out <= 24'h7040a0;
             12'h74b:  out <= 24'h7040b0;
             12'h74c:  out <= 24'h7040c0;
             12'h74d:  out <= 24'h7040d0;
             12'h74e:  out <= 24'h7040e0;
             12'h74f:  out <= 24'h7040f0;
             12'h750:  out <= 24'h705000;
             12'h751:  out <= 24'h705010;
             12'h752:  out <= 24'h705020;
             12'h753:  out <= 24'h705030;
             12'h754:  out <= 24'h705040;
             12'h755:  out <= 24'h705050;
             12'h756:  out <= 24'h705060;
             12'h757:  out <= 24'h705070;
             12'h758:  out <= 24'h705080;
             12'h759:  out <= 24'h705090;
             12'h75a:  out <= 24'h7050a0;
             12'h75b:  out <= 24'h7050b0;
             12'h75c:  out <= 24'h7050c0;
             12'h75d:  out <= 24'h7050d0;
             12'h75e:  out <= 24'h7050e0;
             12'h75f:  out <= 24'h7050f0;
             12'h760:  out <= 24'h706000;
             12'h761:  out <= 24'h706010;
             12'h762:  out <= 24'h706020;
             12'h763:  out <= 24'h706030;
             12'h764:  out <= 24'h706040;
             12'h765:  out <= 24'h706050;
             12'h766:  out <= 24'h706060;
             12'h767:  out <= 24'h706070;
             12'h768:  out <= 24'h706080;
             12'h769:  out <= 24'h706090;
             12'h76a:  out <= 24'h7060a0;
             12'h76b:  out <= 24'h7060b0;
             12'h76c:  out <= 24'h7060c0;
             12'h76d:  out <= 24'h7060d0;
             12'h76e:  out <= 24'h7060e0;
             12'h76f:  out <= 24'h7060f0;
             12'h770:  out <= 24'h707000;
             12'h771:  out <= 24'h707010;
             12'h772:  out <= 24'h707020;
             12'h773:  out <= 24'h707030;
             12'h774:  out <= 24'h707040;
             12'h775:  out <= 24'h707050;
             12'h776:  out <= 24'h707060;
             12'h777:  out <= 24'h707070;
             12'h778:  out <= 24'h707080;
             12'h779:  out <= 24'h707090;
             12'h77a:  out <= 24'h7070a0;
             12'h77b:  out <= 24'h7070b0;
             12'h77c:  out <= 24'h7070c0;
             12'h77d:  out <= 24'h7070d0;
             12'h77e:  out <= 24'h7070e0;
             12'h77f:  out <= 24'h7070f0;
             12'h780:  out <= 24'h708000;
             12'h781:  out <= 24'h708010;
             12'h782:  out <= 24'h708020;
             12'h783:  out <= 24'h708030;
             12'h784:  out <= 24'h708040;
             12'h785:  out <= 24'h708050;
             12'h786:  out <= 24'h708060;
             12'h787:  out <= 24'h708070;
             12'h788:  out <= 24'h708080;
             12'h789:  out <= 24'h708090;
             12'h78a:  out <= 24'h7080a0;
             12'h78b:  out <= 24'h7080b0;
             12'h78c:  out <= 24'h7080c0;
             12'h78d:  out <= 24'h7080d0;
             12'h78e:  out <= 24'h7080e0;
             12'h78f:  out <= 24'h7080f0;
             12'h790:  out <= 24'h709000;
             12'h791:  out <= 24'h709010;
             12'h792:  out <= 24'h709020;
             12'h793:  out <= 24'h709030;
             12'h794:  out <= 24'h709040;
             12'h795:  out <= 24'h709050;
             12'h796:  out <= 24'h709060;
             12'h797:  out <= 24'h709070;
             12'h798:  out <= 24'h709080;
             12'h799:  out <= 24'h709090;
             12'h79a:  out <= 24'h7090a0;
             12'h79b:  out <= 24'h7090b0;
             12'h79c:  out <= 24'h7090c0;
             12'h79d:  out <= 24'h7090d0;
             12'h79e:  out <= 24'h7090e0;
             12'h79f:  out <= 24'h7090f0;
             12'h7a0:  out <= 24'h70a000;
             12'h7a1:  out <= 24'h70a010;
             12'h7a2:  out <= 24'h70a020;
             12'h7a3:  out <= 24'h70a030;
             12'h7a4:  out <= 24'h70a040;
             12'h7a5:  out <= 24'h70a050;
             12'h7a6:  out <= 24'h70a060;
             12'h7a7:  out <= 24'h70a070;
             12'h7a8:  out <= 24'h70a080;
             12'h7a9:  out <= 24'h70a090;
             12'h7aa:  out <= 24'h70a0a0;
             12'h7ab:  out <= 24'h70a0b0;
             12'h7ac:  out <= 24'h70a0c0;
             12'h7ad:  out <= 24'h70a0d0;
             12'h7ae:  out <= 24'h70a0e0;
             12'h7af:  out <= 24'h70a0f0;
             12'h7b0:  out <= 24'h70b000;
             12'h7b1:  out <= 24'h70b010;
             12'h7b2:  out <= 24'h70b020;
             12'h7b3:  out <= 24'h70b030;
             12'h7b4:  out <= 24'h70b040;
             12'h7b5:  out <= 24'h70b050;
             12'h7b6:  out <= 24'h70b060;
             12'h7b7:  out <= 24'h70b070;
             12'h7b8:  out <= 24'h70b080;
             12'h7b9:  out <= 24'h70b090;
             12'h7ba:  out <= 24'h70b0a0;
             12'h7bb:  out <= 24'h70b0b0;
             12'h7bc:  out <= 24'h70b0c0;
             12'h7bd:  out <= 24'h70b0d0;
             12'h7be:  out <= 24'h70b0e0;
             12'h7bf:  out <= 24'h70b0f0;
             12'h7c0:  out <= 24'h70c000;
             12'h7c1:  out <= 24'h70c010;
             12'h7c2:  out <= 24'h70c020;
             12'h7c3:  out <= 24'h70c030;
             12'h7c4:  out <= 24'h70c040;
             12'h7c5:  out <= 24'h70c050;
             12'h7c6:  out <= 24'h70c060;
             12'h7c7:  out <= 24'h70c070;
             12'h7c8:  out <= 24'h70c080;
             12'h7c9:  out <= 24'h70c090;
             12'h7ca:  out <= 24'h70c0a0;
             12'h7cb:  out <= 24'h70c0b0;
             12'h7cc:  out <= 24'h70c0c0;
             12'h7cd:  out <= 24'h70c0d0;
             12'h7ce:  out <= 24'h70c0e0;
             12'h7cf:  out <= 24'h70c0f0;
             12'h7d0:  out <= 24'h70d000;
             12'h7d1:  out <= 24'h70d010;
             12'h7d2:  out <= 24'h70d020;
             12'h7d3:  out <= 24'h70d030;
             12'h7d4:  out <= 24'h70d040;
             12'h7d5:  out <= 24'h70d050;
             12'h7d6:  out <= 24'h70d060;
             12'h7d7:  out <= 24'h70d070;
             12'h7d8:  out <= 24'h70d080;
             12'h7d9:  out <= 24'h70d090;
             12'h7da:  out <= 24'h70d0a0;
             12'h7db:  out <= 24'h70d0b0;
             12'h7dc:  out <= 24'h70d0c0;
             12'h7dd:  out <= 24'h70d0d0;
             12'h7de:  out <= 24'h70d0e0;
             12'h7df:  out <= 24'h70d0f0;
             12'h7e0:  out <= 24'h70e000;
             12'h7e1:  out <= 24'h70e010;
             12'h7e2:  out <= 24'h70e020;
             12'h7e3:  out <= 24'h70e030;
             12'h7e4:  out <= 24'h70e040;
             12'h7e5:  out <= 24'h70e050;
             12'h7e6:  out <= 24'h70e060;
             12'h7e7:  out <= 24'h70e070;
             12'h7e8:  out <= 24'h70e080;
             12'h7e9:  out <= 24'h70e090;
             12'h7ea:  out <= 24'h70e0a0;
             12'h7eb:  out <= 24'h70e0b0;
             12'h7ec:  out <= 24'h70e0c0;
             12'h7ed:  out <= 24'h70e0d0;
             12'h7ee:  out <= 24'h70e0e0;
             12'h7ef:  out <= 24'h70e0f0;
             12'h7f0:  out <= 24'h70f000;
             12'h7f1:  out <= 24'h70f010;
             12'h7f2:  out <= 24'h70f020;
             12'h7f3:  out <= 24'h70f030;
             12'h7f4:  out <= 24'h70f040;
             12'h7f5:  out <= 24'h70f050;
             12'h7f6:  out <= 24'h70f060;
             12'h7f7:  out <= 24'h70f070;
             12'h7f8:  out <= 24'h70f080;
             12'h7f9:  out <= 24'h70f090;
             12'h7fa:  out <= 24'h70f0a0;
             12'h7fb:  out <= 24'h70f0b0;
             12'h7fc:  out <= 24'h70f0c0;
             12'h7fd:  out <= 24'h70f0d0;
             12'h7fe:  out <= 24'h70f0e0;
             12'h7ff:  out <= 24'h70f0f0;
             12'h800:  out <= 24'h800000;
             12'h801:  out <= 24'h800010;
             12'h802:  out <= 24'h800020;
             12'h803:  out <= 24'h800030;
             12'h804:  out <= 24'h800040;
             12'h805:  out <= 24'h800050;
             12'h806:  out <= 24'h800060;
             12'h807:  out <= 24'h800070;
             12'h808:  out <= 24'h800080;
             12'h809:  out <= 24'h800090;
             12'h80a:  out <= 24'h8000a0;
             12'h80b:  out <= 24'h8000b0;
             12'h80c:  out <= 24'h8000c0;
             12'h80d:  out <= 24'h8000d0;
             12'h80e:  out <= 24'h8000e0;
             12'h80f:  out <= 24'h8000f0;
             12'h810:  out <= 24'h801000;
             12'h811:  out <= 24'h801010;
             12'h812:  out <= 24'h801020;
             12'h813:  out <= 24'h801030;
             12'h814:  out <= 24'h801040;
             12'h815:  out <= 24'h801050;
             12'h816:  out <= 24'h801060;
             12'h817:  out <= 24'h801070;
             12'h818:  out <= 24'h801080;
             12'h819:  out <= 24'h801090;
             12'h81a:  out <= 24'h8010a0;
             12'h81b:  out <= 24'h8010b0;
             12'h81c:  out <= 24'h8010c0;
             12'h81d:  out <= 24'h8010d0;
             12'h81e:  out <= 24'h8010e0;
             12'h81f:  out <= 24'h8010f0;
             12'h820:  out <= 24'h802000;
             12'h821:  out <= 24'h802010;
             12'h822:  out <= 24'h802020;
             12'h823:  out <= 24'h802030;
             12'h824:  out <= 24'h802040;
             12'h825:  out <= 24'h802050;
             12'h826:  out <= 24'h802060;
             12'h827:  out <= 24'h802070;
             12'h828:  out <= 24'h802080;
             12'h829:  out <= 24'h802090;
             12'h82a:  out <= 24'h8020a0;
             12'h82b:  out <= 24'h8020b0;
             12'h82c:  out <= 24'h8020c0;
             12'h82d:  out <= 24'h8020d0;
             12'h82e:  out <= 24'h8020e0;
             12'h82f:  out <= 24'h8020f0;
             12'h830:  out <= 24'h803000;
             12'h831:  out <= 24'h803010;
             12'h832:  out <= 24'h803020;
             12'h833:  out <= 24'h803030;
             12'h834:  out <= 24'h803040;
             12'h835:  out <= 24'h803050;
             12'h836:  out <= 24'h803060;
             12'h837:  out <= 24'h803070;
             12'h838:  out <= 24'h803080;
             12'h839:  out <= 24'h803090;
             12'h83a:  out <= 24'h8030a0;
             12'h83b:  out <= 24'h8030b0;
             12'h83c:  out <= 24'h8030c0;
             12'h83d:  out <= 24'h8030d0;
             12'h83e:  out <= 24'h8030e0;
             12'h83f:  out <= 24'h8030f0;
             12'h840:  out <= 24'h804000;
             12'h841:  out <= 24'h804010;
             12'h842:  out <= 24'h804020;
             12'h843:  out <= 24'h804030;
             12'h844:  out <= 24'h804040;
             12'h845:  out <= 24'h804050;
             12'h846:  out <= 24'h804060;
             12'h847:  out <= 24'h804070;
             12'h848:  out <= 24'h804080;
             12'h849:  out <= 24'h804090;
             12'h84a:  out <= 24'h8040a0;
             12'h84b:  out <= 24'h8040b0;
             12'h84c:  out <= 24'h8040c0;
             12'h84d:  out <= 24'h8040d0;
             12'h84e:  out <= 24'h8040e0;
             12'h84f:  out <= 24'h8040f0;
             12'h850:  out <= 24'h805000;
             12'h851:  out <= 24'h805010;
             12'h852:  out <= 24'h805020;
             12'h853:  out <= 24'h805030;
             12'h854:  out <= 24'h805040;
             12'h855:  out <= 24'h805050;
             12'h856:  out <= 24'h805060;
             12'h857:  out <= 24'h805070;
             12'h858:  out <= 24'h805080;
             12'h859:  out <= 24'h805090;
             12'h85a:  out <= 24'h8050a0;
             12'h85b:  out <= 24'h8050b0;
             12'h85c:  out <= 24'h8050c0;
             12'h85d:  out <= 24'h8050d0;
             12'h85e:  out <= 24'h8050e0;
             12'h85f:  out <= 24'h8050f0;
             12'h860:  out <= 24'h806000;
             12'h861:  out <= 24'h806010;
             12'h862:  out <= 24'h806020;
             12'h863:  out <= 24'h806030;
             12'h864:  out <= 24'h806040;
             12'h865:  out <= 24'h806050;
             12'h866:  out <= 24'h806060;
             12'h867:  out <= 24'h806070;
             12'h868:  out <= 24'h806080;
             12'h869:  out <= 24'h806090;
             12'h86a:  out <= 24'h8060a0;
             12'h86b:  out <= 24'h8060b0;
             12'h86c:  out <= 24'h8060c0;
             12'h86d:  out <= 24'h8060d0;
             12'h86e:  out <= 24'h8060e0;
             12'h86f:  out <= 24'h8060f0;
             12'h870:  out <= 24'h807000;
             12'h871:  out <= 24'h807010;
             12'h872:  out <= 24'h807020;
             12'h873:  out <= 24'h807030;
             12'h874:  out <= 24'h807040;
             12'h875:  out <= 24'h807050;
             12'h876:  out <= 24'h807060;
             12'h877:  out <= 24'h807070;
             12'h878:  out <= 24'h807080;
             12'h879:  out <= 24'h807090;
             12'h87a:  out <= 24'h8070a0;
             12'h87b:  out <= 24'h8070b0;
             12'h87c:  out <= 24'h8070c0;
             12'h87d:  out <= 24'h8070d0;
             12'h87e:  out <= 24'h8070e0;
             12'h87f:  out <= 24'h8070f0;
             12'h880:  out <= 24'h808000;
             12'h881:  out <= 24'h808010;
             12'h882:  out <= 24'h808020;
             12'h883:  out <= 24'h808030;
             12'h884:  out <= 24'h808040;
             12'h885:  out <= 24'h808050;
             12'h886:  out <= 24'h808060;
             12'h887:  out <= 24'h808070;
             12'h888:  out <= 24'h808080;
             12'h889:  out <= 24'h808090;
             12'h88a:  out <= 24'h8080a0;
             12'h88b:  out <= 24'h8080b0;
             12'h88c:  out <= 24'h8080c0;
             12'h88d:  out <= 24'h8080d0;
             12'h88e:  out <= 24'h8080e0;
             12'h88f:  out <= 24'h8080f0;
             12'h890:  out <= 24'h809000;
             12'h891:  out <= 24'h809010;
             12'h892:  out <= 24'h809020;
             12'h893:  out <= 24'h809030;
             12'h894:  out <= 24'h809040;
             12'h895:  out <= 24'h809050;
             12'h896:  out <= 24'h809060;
             12'h897:  out <= 24'h809070;
             12'h898:  out <= 24'h809080;
             12'h899:  out <= 24'h809090;
             12'h89a:  out <= 24'h8090a0;
             12'h89b:  out <= 24'h8090b0;
             12'h89c:  out <= 24'h8090c0;
             12'h89d:  out <= 24'h8090d0;
             12'h89e:  out <= 24'h8090e0;
             12'h89f:  out <= 24'h8090f0;
             12'h8a0:  out <= 24'h80a000;
             12'h8a1:  out <= 24'h80a010;
             12'h8a2:  out <= 24'h80a020;
             12'h8a3:  out <= 24'h80a030;
             12'h8a4:  out <= 24'h80a040;
             12'h8a5:  out <= 24'h80a050;
             12'h8a6:  out <= 24'h80a060;
             12'h8a7:  out <= 24'h80a070;
             12'h8a8:  out <= 24'h80a080;
             12'h8a9:  out <= 24'h80a090;
             12'h8aa:  out <= 24'h80a0a0;
             12'h8ab:  out <= 24'h80a0b0;
             12'h8ac:  out <= 24'h80a0c0;
             12'h8ad:  out <= 24'h80a0d0;
             12'h8ae:  out <= 24'h80a0e0;
             12'h8af:  out <= 24'h80a0f0;
             12'h8b0:  out <= 24'h80b000;
             12'h8b1:  out <= 24'h80b010;
             12'h8b2:  out <= 24'h80b020;
             12'h8b3:  out <= 24'h80b030;
             12'h8b4:  out <= 24'h80b040;
             12'h8b5:  out <= 24'h80b050;
             12'h8b6:  out <= 24'h80b060;
             12'h8b7:  out <= 24'h80b070;
             12'h8b8:  out <= 24'h80b080;
             12'h8b9:  out <= 24'h80b090;
             12'h8ba:  out <= 24'h80b0a0;
             12'h8bb:  out <= 24'h80b0b0;
             12'h8bc:  out <= 24'h80b0c0;
             12'h8bd:  out <= 24'h80b0d0;
             12'h8be:  out <= 24'h80b0e0;
             12'h8bf:  out <= 24'h80b0f0;
             12'h8c0:  out <= 24'h80c000;
             12'h8c1:  out <= 24'h80c010;
             12'h8c2:  out <= 24'h80c020;
             12'h8c3:  out <= 24'h80c030;
             12'h8c4:  out <= 24'h80c040;
             12'h8c5:  out <= 24'h80c050;
             12'h8c6:  out <= 24'h80c060;
             12'h8c7:  out <= 24'h80c070;
             12'h8c8:  out <= 24'h80c080;
             12'h8c9:  out <= 24'h80c090;
             12'h8ca:  out <= 24'h80c0a0;
             12'h8cb:  out <= 24'h80c0b0;
             12'h8cc:  out <= 24'h80c0c0;
             12'h8cd:  out <= 24'h80c0d0;
             12'h8ce:  out <= 24'h80c0e0;
             12'h8cf:  out <= 24'h80c0f0;
             12'h8d0:  out <= 24'h80d000;
             12'h8d1:  out <= 24'h80d010;
             12'h8d2:  out <= 24'h80d020;
             12'h8d3:  out <= 24'h80d030;
             12'h8d4:  out <= 24'h80d040;
             12'h8d5:  out <= 24'h80d050;
             12'h8d6:  out <= 24'h80d060;
             12'h8d7:  out <= 24'h80d070;
             12'h8d8:  out <= 24'h80d080;
             12'h8d9:  out <= 24'h80d090;
             12'h8da:  out <= 24'h80d0a0;
             12'h8db:  out <= 24'h80d0b0;
             12'h8dc:  out <= 24'h80d0c0;
             12'h8dd:  out <= 24'h80d0d0;
             12'h8de:  out <= 24'h80d0e0;
             12'h8df:  out <= 24'h80d0f0;
             12'h8e0:  out <= 24'h80e000;
             12'h8e1:  out <= 24'h80e010;
             12'h8e2:  out <= 24'h80e020;
             12'h8e3:  out <= 24'h80e030;
             12'h8e4:  out <= 24'h80e040;
             12'h8e5:  out <= 24'h80e050;
             12'h8e6:  out <= 24'h80e060;
             12'h8e7:  out <= 24'h80e070;
             12'h8e8:  out <= 24'h80e080;
             12'h8e9:  out <= 24'h80e090;
             12'h8ea:  out <= 24'h80e0a0;
             12'h8eb:  out <= 24'h80e0b0;
             12'h8ec:  out <= 24'h80e0c0;
             12'h8ed:  out <= 24'h80e0d0;
             12'h8ee:  out <= 24'h80e0e0;
             12'h8ef:  out <= 24'h80e0f0;
             12'h8f0:  out <= 24'h80f000;
             12'h8f1:  out <= 24'h80f010;
             12'h8f2:  out <= 24'h80f020;
             12'h8f3:  out <= 24'h80f030;
             12'h8f4:  out <= 24'h80f040;
             12'h8f5:  out <= 24'h80f050;
             12'h8f6:  out <= 24'h80f060;
             12'h8f7:  out <= 24'h80f070;
             12'h8f8:  out <= 24'h80f080;
             12'h8f9:  out <= 24'h80f090;
             12'h8fa:  out <= 24'h80f0a0;
             12'h8fb:  out <= 24'h80f0b0;
             12'h8fc:  out <= 24'h80f0c0;
             12'h8fd:  out <= 24'h80f0d0;
             12'h8fe:  out <= 24'h80f0e0;
             12'h8ff:  out <= 24'h80f0f0;
             12'h900:  out <= 24'h900000;
             12'h901:  out <= 24'h900010;
             12'h902:  out <= 24'h900020;
             12'h903:  out <= 24'h900030;
             12'h904:  out <= 24'h900040;
             12'h905:  out <= 24'h900050;
             12'h906:  out <= 24'h900060;
             12'h907:  out <= 24'h900070;
             12'h908:  out <= 24'h900080;
             12'h909:  out <= 24'h900090;
             12'h90a:  out <= 24'h9000a0;
             12'h90b:  out <= 24'h9000b0;
             12'h90c:  out <= 24'h9000c0;
             12'h90d:  out <= 24'h9000d0;
             12'h90e:  out <= 24'h9000e0;
             12'h90f:  out <= 24'h9000f0;
             12'h910:  out <= 24'h901000;
             12'h911:  out <= 24'h901010;
             12'h912:  out <= 24'h901020;
             12'h913:  out <= 24'h901030;
             12'h914:  out <= 24'h901040;
             12'h915:  out <= 24'h901050;
             12'h916:  out <= 24'h901060;
             12'h917:  out <= 24'h901070;
             12'h918:  out <= 24'h901080;
             12'h919:  out <= 24'h901090;
             12'h91a:  out <= 24'h9010a0;
             12'h91b:  out <= 24'h9010b0;
             12'h91c:  out <= 24'h9010c0;
             12'h91d:  out <= 24'h9010d0;
             12'h91e:  out <= 24'h9010e0;
             12'h91f:  out <= 24'h9010f0;
             12'h920:  out <= 24'h902000;
             12'h921:  out <= 24'h902010;
             12'h922:  out <= 24'h902020;
             12'h923:  out <= 24'h902030;
             12'h924:  out <= 24'h902040;
             12'h925:  out <= 24'h902050;
             12'h926:  out <= 24'h902060;
             12'h927:  out <= 24'h902070;
             12'h928:  out <= 24'h902080;
             12'h929:  out <= 24'h902090;
             12'h92a:  out <= 24'h9020a0;
             12'h92b:  out <= 24'h9020b0;
             12'h92c:  out <= 24'h9020c0;
             12'h92d:  out <= 24'h9020d0;
             12'h92e:  out <= 24'h9020e0;
             12'h92f:  out <= 24'h9020f0;
             12'h930:  out <= 24'h903000;
             12'h931:  out <= 24'h903010;
             12'h932:  out <= 24'h903020;
             12'h933:  out <= 24'h903030;
             12'h934:  out <= 24'h903040;
             12'h935:  out <= 24'h903050;
             12'h936:  out <= 24'h903060;
             12'h937:  out <= 24'h903070;
             12'h938:  out <= 24'h903080;
             12'h939:  out <= 24'h903090;
             12'h93a:  out <= 24'h9030a0;
             12'h93b:  out <= 24'h9030b0;
             12'h93c:  out <= 24'h9030c0;
             12'h93d:  out <= 24'h9030d0;
             12'h93e:  out <= 24'h9030e0;
             12'h93f:  out <= 24'h9030f0;
             12'h940:  out <= 24'h904000;
             12'h941:  out <= 24'h904010;
             12'h942:  out <= 24'h904020;
             12'h943:  out <= 24'h904030;
             12'h944:  out <= 24'h904040;
             12'h945:  out <= 24'h904050;
             12'h946:  out <= 24'h904060;
             12'h947:  out <= 24'h904070;
             12'h948:  out <= 24'h904080;
             12'h949:  out <= 24'h904090;
             12'h94a:  out <= 24'h9040a0;
             12'h94b:  out <= 24'h9040b0;
             12'h94c:  out <= 24'h9040c0;
             12'h94d:  out <= 24'h9040d0;
             12'h94e:  out <= 24'h9040e0;
             12'h94f:  out <= 24'h9040f0;
             12'h950:  out <= 24'h905000;
             12'h951:  out <= 24'h905010;
             12'h952:  out <= 24'h905020;
             12'h953:  out <= 24'h905030;
             12'h954:  out <= 24'h905040;
             12'h955:  out <= 24'h905050;
             12'h956:  out <= 24'h905060;
             12'h957:  out <= 24'h905070;
             12'h958:  out <= 24'h905080;
             12'h959:  out <= 24'h905090;
             12'h95a:  out <= 24'h9050a0;
             12'h95b:  out <= 24'h9050b0;
             12'h95c:  out <= 24'h9050c0;
             12'h95d:  out <= 24'h9050d0;
             12'h95e:  out <= 24'h9050e0;
             12'h95f:  out <= 24'h9050f0;
             12'h960:  out <= 24'h906000;
             12'h961:  out <= 24'h906010;
             12'h962:  out <= 24'h906020;
             12'h963:  out <= 24'h906030;
             12'h964:  out <= 24'h906040;
             12'h965:  out <= 24'h906050;
             12'h966:  out <= 24'h906060;
             12'h967:  out <= 24'h906070;
             12'h968:  out <= 24'h906080;
             12'h969:  out <= 24'h906090;
             12'h96a:  out <= 24'h9060a0;
             12'h96b:  out <= 24'h9060b0;
             12'h96c:  out <= 24'h9060c0;
             12'h96d:  out <= 24'h9060d0;
             12'h96e:  out <= 24'h9060e0;
             12'h96f:  out <= 24'h9060f0;
             12'h970:  out <= 24'h907000;
             12'h971:  out <= 24'h907010;
             12'h972:  out <= 24'h907020;
             12'h973:  out <= 24'h907030;
             12'h974:  out <= 24'h907040;
             12'h975:  out <= 24'h907050;
             12'h976:  out <= 24'h907060;
             12'h977:  out <= 24'h907070;
             12'h978:  out <= 24'h907080;
             12'h979:  out <= 24'h907090;
             12'h97a:  out <= 24'h9070a0;
             12'h97b:  out <= 24'h9070b0;
             12'h97c:  out <= 24'h9070c0;
             12'h97d:  out <= 24'h9070d0;
             12'h97e:  out <= 24'h9070e0;
             12'h97f:  out <= 24'h9070f0;
             12'h980:  out <= 24'h908000;
             12'h981:  out <= 24'h908010;
             12'h982:  out <= 24'h908020;
             12'h983:  out <= 24'h908030;
             12'h984:  out <= 24'h908040;
             12'h985:  out <= 24'h908050;
             12'h986:  out <= 24'h908060;
             12'h987:  out <= 24'h908070;
             12'h988:  out <= 24'h908080;
             12'h989:  out <= 24'h908090;
             12'h98a:  out <= 24'h9080a0;
             12'h98b:  out <= 24'h9080b0;
             12'h98c:  out <= 24'h9080c0;
             12'h98d:  out <= 24'h9080d0;
             12'h98e:  out <= 24'h9080e0;
             12'h98f:  out <= 24'h9080f0;
             12'h990:  out <= 24'h909000;
             12'h991:  out <= 24'h909010;
             12'h992:  out <= 24'h909020;
             12'h993:  out <= 24'h909030;
             12'h994:  out <= 24'h909040;
             12'h995:  out <= 24'h909050;
             12'h996:  out <= 24'h909060;
             12'h997:  out <= 24'h909070;
             12'h998:  out <= 24'h909080;
             12'h999:  out <= 24'h909090;
             12'h99a:  out <= 24'h9090a0;
             12'h99b:  out <= 24'h9090b0;
             12'h99c:  out <= 24'h9090c0;
             12'h99d:  out <= 24'h9090d0;
             12'h99e:  out <= 24'h9090e0;
             12'h99f:  out <= 24'h9090f0;
             12'h9a0:  out <= 24'h90a000;
             12'h9a1:  out <= 24'h90a010;
             12'h9a2:  out <= 24'h90a020;
             12'h9a3:  out <= 24'h90a030;
             12'h9a4:  out <= 24'h90a040;
             12'h9a5:  out <= 24'h90a050;
             12'h9a6:  out <= 24'h90a060;
             12'h9a7:  out <= 24'h90a070;
             12'h9a8:  out <= 24'h90a080;
             12'h9a9:  out <= 24'h90a090;
             12'h9aa:  out <= 24'h90a0a0;
             12'h9ab:  out <= 24'h90a0b0;
             12'h9ac:  out <= 24'h90a0c0;
             12'h9ad:  out <= 24'h90a0d0;
             12'h9ae:  out <= 24'h90a0e0;
             12'h9af:  out <= 24'h90a0f0;
             12'h9b0:  out <= 24'h90b000;
             12'h9b1:  out <= 24'h90b010;
             12'h9b2:  out <= 24'h90b020;
             12'h9b3:  out <= 24'h90b030;
             12'h9b4:  out <= 24'h90b040;
             12'h9b5:  out <= 24'h90b050;
             12'h9b6:  out <= 24'h90b060;
             12'h9b7:  out <= 24'h90b070;
             12'h9b8:  out <= 24'h90b080;
             12'h9b9:  out <= 24'h90b090;
             12'h9ba:  out <= 24'h90b0a0;
             12'h9bb:  out <= 24'h90b0b0;
             12'h9bc:  out <= 24'h90b0c0;
             12'h9bd:  out <= 24'h90b0d0;
             12'h9be:  out <= 24'h90b0e0;
             12'h9bf:  out <= 24'h90b0f0;
             12'h9c0:  out <= 24'h90c000;
             12'h9c1:  out <= 24'h90c010;
             12'h9c2:  out <= 24'h90c020;
             12'h9c3:  out <= 24'h90c030;
             12'h9c4:  out <= 24'h90c040;
             12'h9c5:  out <= 24'h90c050;
             12'h9c6:  out <= 24'h90c060;
             12'h9c7:  out <= 24'h90c070;
             12'h9c8:  out <= 24'h90c080;
             12'h9c9:  out <= 24'h90c090;
             12'h9ca:  out <= 24'h90c0a0;
             12'h9cb:  out <= 24'h90c0b0;
             12'h9cc:  out <= 24'h90c0c0;
             12'h9cd:  out <= 24'h90c0d0;
             12'h9ce:  out <= 24'h90c0e0;
             12'h9cf:  out <= 24'h90c0f0;
             12'h9d0:  out <= 24'h90d000;
             12'h9d1:  out <= 24'h90d010;
             12'h9d2:  out <= 24'h90d020;
             12'h9d3:  out <= 24'h90d030;
             12'h9d4:  out <= 24'h90d040;
             12'h9d5:  out <= 24'h90d050;
             12'h9d6:  out <= 24'h90d060;
             12'h9d7:  out <= 24'h90d070;
             12'h9d8:  out <= 24'h90d080;
             12'h9d9:  out <= 24'h90d090;
             12'h9da:  out <= 24'h90d0a0;
             12'h9db:  out <= 24'h90d0b0;
             12'h9dc:  out <= 24'h90d0c0;
             12'h9dd:  out <= 24'h90d0d0;
             12'h9de:  out <= 24'h90d0e0;
             12'h9df:  out <= 24'h90d0f0;
             12'h9e0:  out <= 24'h90e000;
             12'h9e1:  out <= 24'h90e010;
             12'h9e2:  out <= 24'h90e020;
             12'h9e3:  out <= 24'h90e030;
             12'h9e4:  out <= 24'h90e040;
             12'h9e5:  out <= 24'h90e050;
             12'h9e6:  out <= 24'h90e060;
             12'h9e7:  out <= 24'h90e070;
             12'h9e8:  out <= 24'h90e080;
             12'h9e9:  out <= 24'h90e090;
             12'h9ea:  out <= 24'h90e0a0;
             12'h9eb:  out <= 24'h90e0b0;
             12'h9ec:  out <= 24'h90e0c0;
             12'h9ed:  out <= 24'h90e0d0;
             12'h9ee:  out <= 24'h90e0e0;
             12'h9ef:  out <= 24'h90e0f0;
             12'h9f0:  out <= 24'h90f000;
             12'h9f1:  out <= 24'h90f010;
             12'h9f2:  out <= 24'h90f020;
             12'h9f3:  out <= 24'h90f030;
             12'h9f4:  out <= 24'h90f040;
             12'h9f5:  out <= 24'h90f050;
             12'h9f6:  out <= 24'h90f060;
             12'h9f7:  out <= 24'h90f070;
             12'h9f8:  out <= 24'h90f080;
             12'h9f9:  out <= 24'h90f090;
             12'h9fa:  out <= 24'h90f0a0;
             12'h9fb:  out <= 24'h90f0b0;
             12'h9fc:  out <= 24'h90f0c0;
             12'h9fd:  out <= 24'h90f0d0;
             12'h9fe:  out <= 24'h90f0e0;
             12'h9ff:  out <= 24'h90f0f0;
             12'ha00:  out <= 24'ha00000;
             12'ha01:  out <= 24'ha00010;
             12'ha02:  out <= 24'ha00020;
             12'ha03:  out <= 24'ha00030;
             12'ha04:  out <= 24'ha00040;
             12'ha05:  out <= 24'ha00050;
             12'ha06:  out <= 24'ha00060;
             12'ha07:  out <= 24'ha00070;
             12'ha08:  out <= 24'ha00080;
             12'ha09:  out <= 24'ha00090;
             12'ha0a:  out <= 24'ha000a0;
             12'ha0b:  out <= 24'ha000b0;
             12'ha0c:  out <= 24'ha000c0;
             12'ha0d:  out <= 24'ha000d0;
             12'ha0e:  out <= 24'ha000e0;
             12'ha0f:  out <= 24'ha000f0;
             12'ha10:  out <= 24'ha01000;
             12'ha11:  out <= 24'ha01010;
             12'ha12:  out <= 24'ha01020;
             12'ha13:  out <= 24'ha01030;
             12'ha14:  out <= 24'ha01040;
             12'ha15:  out <= 24'ha01050;
             12'ha16:  out <= 24'ha01060;
             12'ha17:  out <= 24'ha01070;
             12'ha18:  out <= 24'ha01080;
             12'ha19:  out <= 24'ha01090;
             12'ha1a:  out <= 24'ha010a0;
             12'ha1b:  out <= 24'ha010b0;
             12'ha1c:  out <= 24'ha010c0;
             12'ha1d:  out <= 24'ha010d0;
             12'ha1e:  out <= 24'ha010e0;
             12'ha1f:  out <= 24'ha010f0;
             12'ha20:  out <= 24'ha02000;
             12'ha21:  out <= 24'ha02010;
             12'ha22:  out <= 24'ha02020;
             12'ha23:  out <= 24'ha02030;
             12'ha24:  out <= 24'ha02040;
             12'ha25:  out <= 24'ha02050;
             12'ha26:  out <= 24'ha02060;
             12'ha27:  out <= 24'ha02070;
             12'ha28:  out <= 24'ha02080;
             12'ha29:  out <= 24'ha02090;
             12'ha2a:  out <= 24'ha020a0;
             12'ha2b:  out <= 24'ha020b0;
             12'ha2c:  out <= 24'ha020c0;
             12'ha2d:  out <= 24'ha020d0;
             12'ha2e:  out <= 24'ha020e0;
             12'ha2f:  out <= 24'ha020f0;
             12'ha30:  out <= 24'ha03000;
             12'ha31:  out <= 24'ha03010;
             12'ha32:  out <= 24'ha03020;
             12'ha33:  out <= 24'ha03030;
             12'ha34:  out <= 24'ha03040;
             12'ha35:  out <= 24'ha03050;
             12'ha36:  out <= 24'ha03060;
             12'ha37:  out <= 24'ha03070;
             12'ha38:  out <= 24'ha03080;
             12'ha39:  out <= 24'ha03090;
             12'ha3a:  out <= 24'ha030a0;
             12'ha3b:  out <= 24'ha030b0;
             12'ha3c:  out <= 24'ha030c0;
             12'ha3d:  out <= 24'ha030d0;
             12'ha3e:  out <= 24'ha030e0;
             12'ha3f:  out <= 24'ha030f0;
             12'ha40:  out <= 24'ha04000;
             12'ha41:  out <= 24'ha04010;
             12'ha42:  out <= 24'ha04020;
             12'ha43:  out <= 24'ha04030;
             12'ha44:  out <= 24'ha04040;
             12'ha45:  out <= 24'ha04050;
             12'ha46:  out <= 24'ha04060;
             12'ha47:  out <= 24'ha04070;
             12'ha48:  out <= 24'ha04080;
             12'ha49:  out <= 24'ha04090;
             12'ha4a:  out <= 24'ha040a0;
             12'ha4b:  out <= 24'ha040b0;
             12'ha4c:  out <= 24'ha040c0;
             12'ha4d:  out <= 24'ha040d0;
             12'ha4e:  out <= 24'ha040e0;
             12'ha4f:  out <= 24'ha040f0;
             12'ha50:  out <= 24'ha05000;
             12'ha51:  out <= 24'ha05010;
             12'ha52:  out <= 24'ha05020;
             12'ha53:  out <= 24'ha05030;
             12'ha54:  out <= 24'ha05040;
             12'ha55:  out <= 24'ha05050;
             12'ha56:  out <= 24'ha05060;
             12'ha57:  out <= 24'ha05070;
             12'ha58:  out <= 24'ha05080;
             12'ha59:  out <= 24'ha05090;
             12'ha5a:  out <= 24'ha050a0;
             12'ha5b:  out <= 24'ha050b0;
             12'ha5c:  out <= 24'ha050c0;
             12'ha5d:  out <= 24'ha050d0;
             12'ha5e:  out <= 24'ha050e0;
             12'ha5f:  out <= 24'ha050f0;
             12'ha60:  out <= 24'ha06000;
             12'ha61:  out <= 24'ha06010;
             12'ha62:  out <= 24'ha06020;
             12'ha63:  out <= 24'ha06030;
             12'ha64:  out <= 24'ha06040;
             12'ha65:  out <= 24'ha06050;
             12'ha66:  out <= 24'ha06060;
             12'ha67:  out <= 24'ha06070;
             12'ha68:  out <= 24'ha06080;
             12'ha69:  out <= 24'ha06090;
             12'ha6a:  out <= 24'ha060a0;
             12'ha6b:  out <= 24'ha060b0;
             12'ha6c:  out <= 24'ha060c0;
             12'ha6d:  out <= 24'ha060d0;
             12'ha6e:  out <= 24'ha060e0;
             12'ha6f:  out <= 24'ha060f0;
             12'ha70:  out <= 24'ha07000;
             12'ha71:  out <= 24'ha07010;
             12'ha72:  out <= 24'ha07020;
             12'ha73:  out <= 24'ha07030;
             12'ha74:  out <= 24'ha07040;
             12'ha75:  out <= 24'ha07050;
             12'ha76:  out <= 24'ha07060;
             12'ha77:  out <= 24'ha07070;
             12'ha78:  out <= 24'ha07080;
             12'ha79:  out <= 24'ha07090;
             12'ha7a:  out <= 24'ha070a0;
             12'ha7b:  out <= 24'ha070b0;
             12'ha7c:  out <= 24'ha070c0;
             12'ha7d:  out <= 24'ha070d0;
             12'ha7e:  out <= 24'ha070e0;
             12'ha7f:  out <= 24'ha070f0;
             12'ha80:  out <= 24'ha08000;
             12'ha81:  out <= 24'ha08010;
             12'ha82:  out <= 24'ha08020;
             12'ha83:  out <= 24'ha08030;
             12'ha84:  out <= 24'ha08040;
             12'ha85:  out <= 24'ha08050;
             12'ha86:  out <= 24'ha08060;
             12'ha87:  out <= 24'ha08070;
             12'ha88:  out <= 24'ha08080;
             12'ha89:  out <= 24'ha08090;
             12'ha8a:  out <= 24'ha080a0;
             12'ha8b:  out <= 24'ha080b0;
             12'ha8c:  out <= 24'ha080c0;
             12'ha8d:  out <= 24'ha080d0;
             12'ha8e:  out <= 24'ha080e0;
             12'ha8f:  out <= 24'ha080f0;
             12'ha90:  out <= 24'ha09000;
             12'ha91:  out <= 24'ha09010;
             12'ha92:  out <= 24'ha09020;
             12'ha93:  out <= 24'ha09030;
             12'ha94:  out <= 24'ha09040;
             12'ha95:  out <= 24'ha09050;
             12'ha96:  out <= 24'ha09060;
             12'ha97:  out <= 24'ha09070;
             12'ha98:  out <= 24'ha09080;
             12'ha99:  out <= 24'ha09090;
             12'ha9a:  out <= 24'ha090a0;
             12'ha9b:  out <= 24'ha090b0;
             12'ha9c:  out <= 24'ha090c0;
             12'ha9d:  out <= 24'ha090d0;
             12'ha9e:  out <= 24'ha090e0;
             12'ha9f:  out <= 24'ha090f0;
             12'haa0:  out <= 24'ha0a000;
             12'haa1:  out <= 24'ha0a010;
             12'haa2:  out <= 24'ha0a020;
             12'haa3:  out <= 24'ha0a030;
             12'haa4:  out <= 24'ha0a040;
             12'haa5:  out <= 24'ha0a050;
             12'haa6:  out <= 24'ha0a060;
             12'haa7:  out <= 24'ha0a070;
             12'haa8:  out <= 24'ha0a080;
             12'haa9:  out <= 24'ha0a090;
             12'haaa:  out <= 24'ha0a0a0;
             12'haab:  out <= 24'ha0a0b0;
             12'haac:  out <= 24'ha0a0c0;
             12'haad:  out <= 24'ha0a0d0;
             12'haae:  out <= 24'ha0a0e0;
             12'haaf:  out <= 24'ha0a0f0;
             12'hab0:  out <= 24'ha0b000;
             12'hab1:  out <= 24'ha0b010;
             12'hab2:  out <= 24'ha0b020;
             12'hab3:  out <= 24'ha0b030;
             12'hab4:  out <= 24'ha0b040;
             12'hab5:  out <= 24'ha0b050;
             12'hab6:  out <= 24'ha0b060;
             12'hab7:  out <= 24'ha0b070;
             12'hab8:  out <= 24'ha0b080;
             12'hab9:  out <= 24'ha0b090;
             12'haba:  out <= 24'ha0b0a0;
             12'habb:  out <= 24'ha0b0b0;
             12'habc:  out <= 24'ha0b0c0;
             12'habd:  out <= 24'ha0b0d0;
             12'habe:  out <= 24'ha0b0e0;
             12'habf:  out <= 24'ha0b0f0;
             12'hac0:  out <= 24'ha0c000;
             12'hac1:  out <= 24'ha0c010;
             12'hac2:  out <= 24'ha0c020;
             12'hac3:  out <= 24'ha0c030;
             12'hac4:  out <= 24'ha0c040;
             12'hac5:  out <= 24'ha0c050;
             12'hac6:  out <= 24'ha0c060;
             12'hac7:  out <= 24'ha0c070;
             12'hac8:  out <= 24'ha0c080;
             12'hac9:  out <= 24'ha0c090;
             12'haca:  out <= 24'ha0c0a0;
             12'hacb:  out <= 24'ha0c0b0;
             12'hacc:  out <= 24'ha0c0c0;
             12'hacd:  out <= 24'ha0c0d0;
             12'hace:  out <= 24'ha0c0e0;
             12'hacf:  out <= 24'ha0c0f0;
             12'had0:  out <= 24'ha0d000;
             12'had1:  out <= 24'ha0d010;
             12'had2:  out <= 24'ha0d020;
             12'had3:  out <= 24'ha0d030;
             12'had4:  out <= 24'ha0d040;
             12'had5:  out <= 24'ha0d050;
             12'had6:  out <= 24'ha0d060;
             12'had7:  out <= 24'ha0d070;
             12'had8:  out <= 24'ha0d080;
             12'had9:  out <= 24'ha0d090;
             12'hada:  out <= 24'ha0d0a0;
             12'hadb:  out <= 24'ha0d0b0;
             12'hadc:  out <= 24'ha0d0c0;
             12'hadd:  out <= 24'ha0d0d0;
             12'hade:  out <= 24'ha0d0e0;
             12'hadf:  out <= 24'ha0d0f0;
             12'hae0:  out <= 24'ha0e000;
             12'hae1:  out <= 24'ha0e010;
             12'hae2:  out <= 24'ha0e020;
             12'hae3:  out <= 24'ha0e030;
             12'hae4:  out <= 24'ha0e040;
             12'hae5:  out <= 24'ha0e050;
             12'hae6:  out <= 24'ha0e060;
             12'hae7:  out <= 24'ha0e070;
             12'hae8:  out <= 24'ha0e080;
             12'hae9:  out <= 24'ha0e090;
             12'haea:  out <= 24'ha0e0a0;
             12'haeb:  out <= 24'ha0e0b0;
             12'haec:  out <= 24'ha0e0c0;
             12'haed:  out <= 24'ha0e0d0;
             12'haee:  out <= 24'ha0e0e0;
             12'haef:  out <= 24'ha0e0f0;
             12'haf0:  out <= 24'ha0f000;
             12'haf1:  out <= 24'ha0f010;
             12'haf2:  out <= 24'ha0f020;
             12'haf3:  out <= 24'ha0f030;
             12'haf4:  out <= 24'ha0f040;
             12'haf5:  out <= 24'ha0f050;
             12'haf6:  out <= 24'ha0f060;
             12'haf7:  out <= 24'ha0f070;
             12'haf8:  out <= 24'ha0f080;
             12'haf9:  out <= 24'ha0f090;
             12'hafa:  out <= 24'ha0f0a0;
             12'hafb:  out <= 24'ha0f0b0;
             12'hafc:  out <= 24'ha0f0c0;
             12'hafd:  out <= 24'ha0f0d0;
             12'hafe:  out <= 24'ha0f0e0;
             12'haff:  out <= 24'ha0f0f0;
             12'hb00:  out <= 24'hb00000;
             12'hb01:  out <= 24'hb00010;
             12'hb02:  out <= 24'hb00020;
             12'hb03:  out <= 24'hb00030;
             12'hb04:  out <= 24'hb00040;
             12'hb05:  out <= 24'hb00050;
             12'hb06:  out <= 24'hb00060;
             12'hb07:  out <= 24'hb00070;
             12'hb08:  out <= 24'hb00080;
             12'hb09:  out <= 24'hb00090;
             12'hb0a:  out <= 24'hb000a0;
             12'hb0b:  out <= 24'hb000b0;
             12'hb0c:  out <= 24'hb000c0;
             12'hb0d:  out <= 24'hb000d0;
             12'hb0e:  out <= 24'hb000e0;
             12'hb0f:  out <= 24'hb000f0;
             12'hb10:  out <= 24'hb01000;
             12'hb11:  out <= 24'hb01010;
             12'hb12:  out <= 24'hb01020;
             12'hb13:  out <= 24'hb01030;
             12'hb14:  out <= 24'hb01040;
             12'hb15:  out <= 24'hb01050;
             12'hb16:  out <= 24'hb01060;
             12'hb17:  out <= 24'hb01070;
             12'hb18:  out <= 24'hb01080;
             12'hb19:  out <= 24'hb01090;
             12'hb1a:  out <= 24'hb010a0;
             12'hb1b:  out <= 24'hb010b0;
             12'hb1c:  out <= 24'hb010c0;
             12'hb1d:  out <= 24'hb010d0;
             12'hb1e:  out <= 24'hb010e0;
             12'hb1f:  out <= 24'hb010f0;
             12'hb20:  out <= 24'hb02000;
             12'hb21:  out <= 24'hb02010;
             12'hb22:  out <= 24'hb02020;
             12'hb23:  out <= 24'hb02030;
             12'hb24:  out <= 24'hb02040;
             12'hb25:  out <= 24'hb02050;
             12'hb26:  out <= 24'hb02060;
             12'hb27:  out <= 24'hb02070;
             12'hb28:  out <= 24'hb02080;
             12'hb29:  out <= 24'hb02090;
             12'hb2a:  out <= 24'hb020a0;
             12'hb2b:  out <= 24'hb020b0;
             12'hb2c:  out <= 24'hb020c0;
             12'hb2d:  out <= 24'hb020d0;
             12'hb2e:  out <= 24'hb020e0;
             12'hb2f:  out <= 24'hb020f0;
             12'hb30:  out <= 24'hb03000;
             12'hb31:  out <= 24'hb03010;
             12'hb32:  out <= 24'hb03020;
             12'hb33:  out <= 24'hb03030;
             12'hb34:  out <= 24'hb03040;
             12'hb35:  out <= 24'hb03050;
             12'hb36:  out <= 24'hb03060;
             12'hb37:  out <= 24'hb03070;
             12'hb38:  out <= 24'hb03080;
             12'hb39:  out <= 24'hb03090;
             12'hb3a:  out <= 24'hb030a0;
             12'hb3b:  out <= 24'hb030b0;
             12'hb3c:  out <= 24'hb030c0;
             12'hb3d:  out <= 24'hb030d0;
             12'hb3e:  out <= 24'hb030e0;
             12'hb3f:  out <= 24'hb030f0;
             12'hb40:  out <= 24'hb04000;
             12'hb41:  out <= 24'hb04010;
             12'hb42:  out <= 24'hb04020;
             12'hb43:  out <= 24'hb04030;
             12'hb44:  out <= 24'hb04040;
             12'hb45:  out <= 24'hb04050;
             12'hb46:  out <= 24'hb04060;
             12'hb47:  out <= 24'hb04070;
             12'hb48:  out <= 24'hb04080;
             12'hb49:  out <= 24'hb04090;
             12'hb4a:  out <= 24'hb040a0;
             12'hb4b:  out <= 24'hb040b0;
             12'hb4c:  out <= 24'hb040c0;
             12'hb4d:  out <= 24'hb040d0;
             12'hb4e:  out <= 24'hb040e0;
             12'hb4f:  out <= 24'hb040f0;
             12'hb50:  out <= 24'hb05000;
             12'hb51:  out <= 24'hb05010;
             12'hb52:  out <= 24'hb05020;
             12'hb53:  out <= 24'hb05030;
             12'hb54:  out <= 24'hb05040;
             12'hb55:  out <= 24'hb05050;
             12'hb56:  out <= 24'hb05060;
             12'hb57:  out <= 24'hb05070;
             12'hb58:  out <= 24'hb05080;
             12'hb59:  out <= 24'hb05090;
             12'hb5a:  out <= 24'hb050a0;
             12'hb5b:  out <= 24'hb050b0;
             12'hb5c:  out <= 24'hb050c0;
             12'hb5d:  out <= 24'hb050d0;
             12'hb5e:  out <= 24'hb050e0;
             12'hb5f:  out <= 24'hb050f0;
             12'hb60:  out <= 24'hb06000;
             12'hb61:  out <= 24'hb06010;
             12'hb62:  out <= 24'hb06020;
             12'hb63:  out <= 24'hb06030;
             12'hb64:  out <= 24'hb06040;
             12'hb65:  out <= 24'hb06050;
             12'hb66:  out <= 24'hb06060;
             12'hb67:  out <= 24'hb06070;
             12'hb68:  out <= 24'hb06080;
             12'hb69:  out <= 24'hb06090;
             12'hb6a:  out <= 24'hb060a0;
             12'hb6b:  out <= 24'hb060b0;
             12'hb6c:  out <= 24'hb060c0;
             12'hb6d:  out <= 24'hb060d0;
             12'hb6e:  out <= 24'hb060e0;
             12'hb6f:  out <= 24'hb060f0;
             12'hb70:  out <= 24'hb07000;
             12'hb71:  out <= 24'hb07010;
             12'hb72:  out <= 24'hb07020;
             12'hb73:  out <= 24'hb07030;
             12'hb74:  out <= 24'hb07040;
             12'hb75:  out <= 24'hb07050;
             12'hb76:  out <= 24'hb07060;
             12'hb77:  out <= 24'hb07070;
             12'hb78:  out <= 24'hb07080;
             12'hb79:  out <= 24'hb07090;
             12'hb7a:  out <= 24'hb070a0;
             12'hb7b:  out <= 24'hb070b0;
             12'hb7c:  out <= 24'hb070c0;
             12'hb7d:  out <= 24'hb070d0;
             12'hb7e:  out <= 24'hb070e0;
             12'hb7f:  out <= 24'hb070f0;
             12'hb80:  out <= 24'hb08000;
             12'hb81:  out <= 24'hb08010;
             12'hb82:  out <= 24'hb08020;
             12'hb83:  out <= 24'hb08030;
             12'hb84:  out <= 24'hb08040;
             12'hb85:  out <= 24'hb08050;
             12'hb86:  out <= 24'hb08060;
             12'hb87:  out <= 24'hb08070;
             12'hb88:  out <= 24'hb08080;
             12'hb89:  out <= 24'hb08090;
             12'hb8a:  out <= 24'hb080a0;
             12'hb8b:  out <= 24'hb080b0;
             12'hb8c:  out <= 24'hb080c0;
             12'hb8d:  out <= 24'hb080d0;
             12'hb8e:  out <= 24'hb080e0;
             12'hb8f:  out <= 24'hb080f0;
             12'hb90:  out <= 24'hb09000;
             12'hb91:  out <= 24'hb09010;
             12'hb92:  out <= 24'hb09020;
             12'hb93:  out <= 24'hb09030;
             12'hb94:  out <= 24'hb09040;
             12'hb95:  out <= 24'hb09050;
             12'hb96:  out <= 24'hb09060;
             12'hb97:  out <= 24'hb09070;
             12'hb98:  out <= 24'hb09080;
             12'hb99:  out <= 24'hb09090;
             12'hb9a:  out <= 24'hb090a0;
             12'hb9b:  out <= 24'hb090b0;
             12'hb9c:  out <= 24'hb090c0;
             12'hb9d:  out <= 24'hb090d0;
             12'hb9e:  out <= 24'hb090e0;
             12'hb9f:  out <= 24'hb090f0;
             12'hba0:  out <= 24'hb0a000;
             12'hba1:  out <= 24'hb0a010;
             12'hba2:  out <= 24'hb0a020;
             12'hba3:  out <= 24'hb0a030;
             12'hba4:  out <= 24'hb0a040;
             12'hba5:  out <= 24'hb0a050;
             12'hba6:  out <= 24'hb0a060;
             12'hba7:  out <= 24'hb0a070;
             12'hba8:  out <= 24'hb0a080;
             12'hba9:  out <= 24'hb0a090;
             12'hbaa:  out <= 24'hb0a0a0;
             12'hbab:  out <= 24'hb0a0b0;
             12'hbac:  out <= 24'hb0a0c0;
             12'hbad:  out <= 24'hb0a0d0;
             12'hbae:  out <= 24'hb0a0e0;
             12'hbaf:  out <= 24'hb0a0f0;
             12'hbb0:  out <= 24'hb0b000;
             12'hbb1:  out <= 24'hb0b010;
             12'hbb2:  out <= 24'hb0b020;
             12'hbb3:  out <= 24'hb0b030;
             12'hbb4:  out <= 24'hb0b040;
             12'hbb5:  out <= 24'hb0b050;
             12'hbb6:  out <= 24'hb0b060;
             12'hbb7:  out <= 24'hb0b070;
             12'hbb8:  out <= 24'hb0b080;
             12'hbb9:  out <= 24'hb0b090;
             12'hbba:  out <= 24'hb0b0a0;
             12'hbbb:  out <= 24'hb0b0b0;
             12'hbbc:  out <= 24'hb0b0c0;
             12'hbbd:  out <= 24'hb0b0d0;
             12'hbbe:  out <= 24'hb0b0e0;
             12'hbbf:  out <= 24'hb0b0f0;
             12'hbc0:  out <= 24'hb0c000;
             12'hbc1:  out <= 24'hb0c010;
             12'hbc2:  out <= 24'hb0c020;
             12'hbc3:  out <= 24'hb0c030;
             12'hbc4:  out <= 24'hb0c040;
             12'hbc5:  out <= 24'hb0c050;
             12'hbc6:  out <= 24'hb0c060;
             12'hbc7:  out <= 24'hb0c070;
             12'hbc8:  out <= 24'hb0c080;
             12'hbc9:  out <= 24'hb0c090;
             12'hbca:  out <= 24'hb0c0a0;
             12'hbcb:  out <= 24'hb0c0b0;
             12'hbcc:  out <= 24'hb0c0c0;
             12'hbcd:  out <= 24'hb0c0d0;
             12'hbce:  out <= 24'hb0c0e0;
             12'hbcf:  out <= 24'hb0c0f0;
             12'hbd0:  out <= 24'hb0d000;
             12'hbd1:  out <= 24'hb0d010;
             12'hbd2:  out <= 24'hb0d020;
             12'hbd3:  out <= 24'hb0d030;
             12'hbd4:  out <= 24'hb0d040;
             12'hbd5:  out <= 24'hb0d050;
             12'hbd6:  out <= 24'hb0d060;
             12'hbd7:  out <= 24'hb0d070;
             12'hbd8:  out <= 24'hb0d080;
             12'hbd9:  out <= 24'hb0d090;
             12'hbda:  out <= 24'hb0d0a0;
             12'hbdb:  out <= 24'hb0d0b0;
             12'hbdc:  out <= 24'hb0d0c0;
             12'hbdd:  out <= 24'hb0d0d0;
             12'hbde:  out <= 24'hb0d0e0;
             12'hbdf:  out <= 24'hb0d0f0;
             12'hbe0:  out <= 24'hb0e000;
             12'hbe1:  out <= 24'hb0e010;
             12'hbe2:  out <= 24'hb0e020;
             12'hbe3:  out <= 24'hb0e030;
             12'hbe4:  out <= 24'hb0e040;
             12'hbe5:  out <= 24'hb0e050;
             12'hbe6:  out <= 24'hb0e060;
             12'hbe7:  out <= 24'hb0e070;
             12'hbe8:  out <= 24'hb0e080;
             12'hbe9:  out <= 24'hb0e090;
             12'hbea:  out <= 24'hb0e0a0;
             12'hbeb:  out <= 24'hb0e0b0;
             12'hbec:  out <= 24'hb0e0c0;
             12'hbed:  out <= 24'hb0e0d0;
             12'hbee:  out <= 24'hb0e0e0;
             12'hbef:  out <= 24'hb0e0f0;
             12'hbf0:  out <= 24'hb0f000;
             12'hbf1:  out <= 24'hb0f010;
             12'hbf2:  out <= 24'hb0f020;
             12'hbf3:  out <= 24'hb0f030;
             12'hbf4:  out <= 24'hb0f040;
             12'hbf5:  out <= 24'hb0f050;
             12'hbf6:  out <= 24'hb0f060;
             12'hbf7:  out <= 24'hb0f070;
             12'hbf8:  out <= 24'hb0f080;
             12'hbf9:  out <= 24'hb0f090;
             12'hbfa:  out <= 24'hb0f0a0;
             12'hbfb:  out <= 24'hb0f0b0;
             12'hbfc:  out <= 24'hb0f0c0;
             12'hbfd:  out <= 24'hb0f0d0;
             12'hbfe:  out <= 24'hb0f0e0;
             12'hbff:  out <= 24'hb0f0f0;
             12'hc00:  out <= 24'hc00000;
             12'hc01:  out <= 24'hc00010;
             12'hc02:  out <= 24'hc00020;
             12'hc03:  out <= 24'hc00030;
             12'hc04:  out <= 24'hc00040;
             12'hc05:  out <= 24'hc00050;
             12'hc06:  out <= 24'hc00060;
             12'hc07:  out <= 24'hc00070;
             12'hc08:  out <= 24'hc00080;
             12'hc09:  out <= 24'hc00090;
             12'hc0a:  out <= 24'hc000a0;
             12'hc0b:  out <= 24'hc000b0;
             12'hc0c:  out <= 24'hc000c0;
             12'hc0d:  out <= 24'hc000d0;
             12'hc0e:  out <= 24'hc000e0;
             12'hc0f:  out <= 24'hc000f0;
             12'hc10:  out <= 24'hc01000;
             12'hc11:  out <= 24'hc01010;
             12'hc12:  out <= 24'hc01020;
             12'hc13:  out <= 24'hc01030;
             12'hc14:  out <= 24'hc01040;
             12'hc15:  out <= 24'hc01050;
             12'hc16:  out <= 24'hc01060;
             12'hc17:  out <= 24'hc01070;
             12'hc18:  out <= 24'hc01080;
             12'hc19:  out <= 24'hc01090;
             12'hc1a:  out <= 24'hc010a0;
             12'hc1b:  out <= 24'hc010b0;
             12'hc1c:  out <= 24'hc010c0;
             12'hc1d:  out <= 24'hc010d0;
             12'hc1e:  out <= 24'hc010e0;
             12'hc1f:  out <= 24'hc010f0;
             12'hc20:  out <= 24'hc02000;
             12'hc21:  out <= 24'hc02010;
             12'hc22:  out <= 24'hc02020;
             12'hc23:  out <= 24'hc02030;
             12'hc24:  out <= 24'hc02040;
             12'hc25:  out <= 24'hc02050;
             12'hc26:  out <= 24'hc02060;
             12'hc27:  out <= 24'hc02070;
             12'hc28:  out <= 24'hc02080;
             12'hc29:  out <= 24'hc02090;
             12'hc2a:  out <= 24'hc020a0;
             12'hc2b:  out <= 24'hc020b0;
             12'hc2c:  out <= 24'hc020c0;
             12'hc2d:  out <= 24'hc020d0;
             12'hc2e:  out <= 24'hc020e0;
             12'hc2f:  out <= 24'hc020f0;
             12'hc30:  out <= 24'hc03000;
             12'hc31:  out <= 24'hc03010;
             12'hc32:  out <= 24'hc03020;
             12'hc33:  out <= 24'hc03030;
             12'hc34:  out <= 24'hc03040;
             12'hc35:  out <= 24'hc03050;
             12'hc36:  out <= 24'hc03060;
             12'hc37:  out <= 24'hc03070;
             12'hc38:  out <= 24'hc03080;
             12'hc39:  out <= 24'hc03090;
             12'hc3a:  out <= 24'hc030a0;
             12'hc3b:  out <= 24'hc030b0;
             12'hc3c:  out <= 24'hc030c0;
             12'hc3d:  out <= 24'hc030d0;
             12'hc3e:  out <= 24'hc030e0;
             12'hc3f:  out <= 24'hc030f0;
             12'hc40:  out <= 24'hc04000;
             12'hc41:  out <= 24'hc04010;
             12'hc42:  out <= 24'hc04020;
             12'hc43:  out <= 24'hc04030;
             12'hc44:  out <= 24'hc04040;
             12'hc45:  out <= 24'hc04050;
             12'hc46:  out <= 24'hc04060;
             12'hc47:  out <= 24'hc04070;
             12'hc48:  out <= 24'hc04080;
             12'hc49:  out <= 24'hc04090;
             12'hc4a:  out <= 24'hc040a0;
             12'hc4b:  out <= 24'hc040b0;
             12'hc4c:  out <= 24'hc040c0;
             12'hc4d:  out <= 24'hc040d0;
             12'hc4e:  out <= 24'hc040e0;
             12'hc4f:  out <= 24'hc040f0;
             12'hc50:  out <= 24'hc05000;
             12'hc51:  out <= 24'hc05010;
             12'hc52:  out <= 24'hc05020;
             12'hc53:  out <= 24'hc05030;
             12'hc54:  out <= 24'hc05040;
             12'hc55:  out <= 24'hc05050;
             12'hc56:  out <= 24'hc05060;
             12'hc57:  out <= 24'hc05070;
             12'hc58:  out <= 24'hc05080;
             12'hc59:  out <= 24'hc05090;
             12'hc5a:  out <= 24'hc050a0;
             12'hc5b:  out <= 24'hc050b0;
             12'hc5c:  out <= 24'hc050c0;
             12'hc5d:  out <= 24'hc050d0;
             12'hc5e:  out <= 24'hc050e0;
             12'hc5f:  out <= 24'hc050f0;
             12'hc60:  out <= 24'hc06000;
             12'hc61:  out <= 24'hc06010;
             12'hc62:  out <= 24'hc06020;
             12'hc63:  out <= 24'hc06030;
             12'hc64:  out <= 24'hc06040;
             12'hc65:  out <= 24'hc06050;
             12'hc66:  out <= 24'hc06060;
             12'hc67:  out <= 24'hc06070;
             12'hc68:  out <= 24'hc06080;
             12'hc69:  out <= 24'hc06090;
             12'hc6a:  out <= 24'hc060a0;
             12'hc6b:  out <= 24'hc060b0;
             12'hc6c:  out <= 24'hc060c0;
             12'hc6d:  out <= 24'hc060d0;
             12'hc6e:  out <= 24'hc060e0;
             12'hc6f:  out <= 24'hc060f0;
             12'hc70:  out <= 24'hc07000;
             12'hc71:  out <= 24'hc07010;
             12'hc72:  out <= 24'hc07020;
             12'hc73:  out <= 24'hc07030;
             12'hc74:  out <= 24'hc07040;
             12'hc75:  out <= 24'hc07050;
             12'hc76:  out <= 24'hc07060;
             12'hc77:  out <= 24'hc07070;
             12'hc78:  out <= 24'hc07080;
             12'hc79:  out <= 24'hc07090;
             12'hc7a:  out <= 24'hc070a0;
             12'hc7b:  out <= 24'hc070b0;
             12'hc7c:  out <= 24'hc070c0;
             12'hc7d:  out <= 24'hc070d0;
             12'hc7e:  out <= 24'hc070e0;
             12'hc7f:  out <= 24'hc070f0;
             12'hc80:  out <= 24'hc08000;
             12'hc81:  out <= 24'hc08010;
             12'hc82:  out <= 24'hc08020;
             12'hc83:  out <= 24'hc08030;
             12'hc84:  out <= 24'hc08040;
             12'hc85:  out <= 24'hc08050;
             12'hc86:  out <= 24'hc08060;
             12'hc87:  out <= 24'hc08070;
             12'hc88:  out <= 24'hc08080;
             12'hc89:  out <= 24'hc08090;
             12'hc8a:  out <= 24'hc080a0;
             12'hc8b:  out <= 24'hc080b0;
             12'hc8c:  out <= 24'hc080c0;
             12'hc8d:  out <= 24'hc080d0;
             12'hc8e:  out <= 24'hc080e0;
             12'hc8f:  out <= 24'hc080f0;
             12'hc90:  out <= 24'hc09000;
             12'hc91:  out <= 24'hc09010;
             12'hc92:  out <= 24'hc09020;
             12'hc93:  out <= 24'hc09030;
             12'hc94:  out <= 24'hc09040;
             12'hc95:  out <= 24'hc09050;
             12'hc96:  out <= 24'hc09060;
             12'hc97:  out <= 24'hc09070;
             12'hc98:  out <= 24'hc09080;
             12'hc99:  out <= 24'hc09090;
             12'hc9a:  out <= 24'hc090a0;
             12'hc9b:  out <= 24'hc090b0;
             12'hc9c:  out <= 24'hc090c0;
             12'hc9d:  out <= 24'hc090d0;
             12'hc9e:  out <= 24'hc090e0;
             12'hc9f:  out <= 24'hc090f0;
             12'hca0:  out <= 24'hc0a000;
             12'hca1:  out <= 24'hc0a010;
             12'hca2:  out <= 24'hc0a020;
             12'hca3:  out <= 24'hc0a030;
             12'hca4:  out <= 24'hc0a040;
             12'hca5:  out <= 24'hc0a050;
             12'hca6:  out <= 24'hc0a060;
             12'hca7:  out <= 24'hc0a070;
             12'hca8:  out <= 24'hc0a080;
             12'hca9:  out <= 24'hc0a090;
             12'hcaa:  out <= 24'hc0a0a0;
             12'hcab:  out <= 24'hc0a0b0;
             12'hcac:  out <= 24'hc0a0c0;
             12'hcad:  out <= 24'hc0a0d0;
             12'hcae:  out <= 24'hc0a0e0;
             12'hcaf:  out <= 24'hc0a0f0;
             12'hcb0:  out <= 24'hc0b000;
             12'hcb1:  out <= 24'hc0b010;
             12'hcb2:  out <= 24'hc0b020;
             12'hcb3:  out <= 24'hc0b030;
             12'hcb4:  out <= 24'hc0b040;
             12'hcb5:  out <= 24'hc0b050;
             12'hcb6:  out <= 24'hc0b060;
             12'hcb7:  out <= 24'hc0b070;
             12'hcb8:  out <= 24'hc0b080;
             12'hcb9:  out <= 24'hc0b090;
             12'hcba:  out <= 24'hc0b0a0;
             12'hcbb:  out <= 24'hc0b0b0;
             12'hcbc:  out <= 24'hc0b0c0;
             12'hcbd:  out <= 24'hc0b0d0;
             12'hcbe:  out <= 24'hc0b0e0;
             12'hcbf:  out <= 24'hc0b0f0;
             12'hcc0:  out <= 24'hc0c000;
             12'hcc1:  out <= 24'hc0c010;
             12'hcc2:  out <= 24'hc0c020;
             12'hcc3:  out <= 24'hc0c030;
             12'hcc4:  out <= 24'hc0c040;
             12'hcc5:  out <= 24'hc0c050;
             12'hcc6:  out <= 24'hc0c060;
             12'hcc7:  out <= 24'hc0c070;
             12'hcc8:  out <= 24'hc0c080;
             12'hcc9:  out <= 24'hc0c090;
             12'hcca:  out <= 24'hc0c0a0;
             12'hccb:  out <= 24'hc0c0b0;
             12'hccc:  out <= 24'hc0c0c0;
             12'hccd:  out <= 24'hc0c0d0;
             12'hcce:  out <= 24'hc0c0e0;
             12'hccf:  out <= 24'hc0c0f0;
             12'hcd0:  out <= 24'hc0d000;
             12'hcd1:  out <= 24'hc0d010;
             12'hcd2:  out <= 24'hc0d020;
             12'hcd3:  out <= 24'hc0d030;
             12'hcd4:  out <= 24'hc0d040;
             12'hcd5:  out <= 24'hc0d050;
             12'hcd6:  out <= 24'hc0d060;
             12'hcd7:  out <= 24'hc0d070;
             12'hcd8:  out <= 24'hc0d080;
             12'hcd9:  out <= 24'hc0d090;
             12'hcda:  out <= 24'hc0d0a0;
             12'hcdb:  out <= 24'hc0d0b0;
             12'hcdc:  out <= 24'hc0d0c0;
             12'hcdd:  out <= 24'hc0d0d0;
             12'hcde:  out <= 24'hc0d0e0;
             12'hcdf:  out <= 24'hc0d0f0;
             12'hce0:  out <= 24'hc0e000;
             12'hce1:  out <= 24'hc0e010;
             12'hce2:  out <= 24'hc0e020;
             12'hce3:  out <= 24'hc0e030;
             12'hce4:  out <= 24'hc0e040;
             12'hce5:  out <= 24'hc0e050;
             12'hce6:  out <= 24'hc0e060;
             12'hce7:  out <= 24'hc0e070;
             12'hce8:  out <= 24'hc0e080;
             12'hce9:  out <= 24'hc0e090;
             12'hcea:  out <= 24'hc0e0a0;
             12'hceb:  out <= 24'hc0e0b0;
             12'hcec:  out <= 24'hc0e0c0;
             12'hced:  out <= 24'hc0e0d0;
             12'hcee:  out <= 24'hc0e0e0;
             12'hcef:  out <= 24'hc0e0f0;
             12'hcf0:  out <= 24'hc0f000;
             12'hcf1:  out <= 24'hc0f010;
             12'hcf2:  out <= 24'hc0f020;
             12'hcf3:  out <= 24'hc0f030;
             12'hcf4:  out <= 24'hc0f040;
             12'hcf5:  out <= 24'hc0f050;
             12'hcf6:  out <= 24'hc0f060;
             12'hcf7:  out <= 24'hc0f070;
             12'hcf8:  out <= 24'hc0f080;
             12'hcf9:  out <= 24'hc0f090;
             12'hcfa:  out <= 24'hc0f0a0;
             12'hcfb:  out <= 24'hc0f0b0;
             12'hcfc:  out <= 24'hc0f0c0;
             12'hcfd:  out <= 24'hc0f0d0;
             12'hcfe:  out <= 24'hc0f0e0;
             12'hcff:  out <= 24'hc0f0f0;
             12'hd00:  out <= 24'hd00000;
             12'hd01:  out <= 24'hd00010;
             12'hd02:  out <= 24'hd00020;
             12'hd03:  out <= 24'hd00030;
             12'hd04:  out <= 24'hd00040;
             12'hd05:  out <= 24'hd00050;
             12'hd06:  out <= 24'hd00060;
             12'hd07:  out <= 24'hd00070;
             12'hd08:  out <= 24'hd00080;
             12'hd09:  out <= 24'hd00090;
             12'hd0a:  out <= 24'hd000a0;
             12'hd0b:  out <= 24'hd000b0;
             12'hd0c:  out <= 24'hd000c0;
             12'hd0d:  out <= 24'hd000d0;
             12'hd0e:  out <= 24'hd000e0;
             12'hd0f:  out <= 24'hd000f0;
             12'hd10:  out <= 24'hd01000;
             12'hd11:  out <= 24'hd01010;
             12'hd12:  out <= 24'hd01020;
             12'hd13:  out <= 24'hd01030;
             12'hd14:  out <= 24'hd01040;
             12'hd15:  out <= 24'hd01050;
             12'hd16:  out <= 24'hd01060;
             12'hd17:  out <= 24'hd01070;
             12'hd18:  out <= 24'hd01080;
             12'hd19:  out <= 24'hd01090;
             12'hd1a:  out <= 24'hd010a0;
             12'hd1b:  out <= 24'hd010b0;
             12'hd1c:  out <= 24'hd010c0;
             12'hd1d:  out <= 24'hd010d0;
             12'hd1e:  out <= 24'hd010e0;
             12'hd1f:  out <= 24'hd010f0;
             12'hd20:  out <= 24'hd02000;
             12'hd21:  out <= 24'hd02010;
             12'hd22:  out <= 24'hd02020;
             12'hd23:  out <= 24'hd02030;
             12'hd24:  out <= 24'hd02040;
             12'hd25:  out <= 24'hd02050;
             12'hd26:  out <= 24'hd02060;
             12'hd27:  out <= 24'hd02070;
             12'hd28:  out <= 24'hd02080;
             12'hd29:  out <= 24'hd02090;
             12'hd2a:  out <= 24'hd020a0;
             12'hd2b:  out <= 24'hd020b0;
             12'hd2c:  out <= 24'hd020c0;
             12'hd2d:  out <= 24'hd020d0;
             12'hd2e:  out <= 24'hd020e0;
             12'hd2f:  out <= 24'hd020f0;
             12'hd30:  out <= 24'hd03000;
             12'hd31:  out <= 24'hd03010;
             12'hd32:  out <= 24'hd03020;
             12'hd33:  out <= 24'hd03030;
             12'hd34:  out <= 24'hd03040;
             12'hd35:  out <= 24'hd03050;
             12'hd36:  out <= 24'hd03060;
             12'hd37:  out <= 24'hd03070;
             12'hd38:  out <= 24'hd03080;
             12'hd39:  out <= 24'hd03090;
             12'hd3a:  out <= 24'hd030a0;
             12'hd3b:  out <= 24'hd030b0;
             12'hd3c:  out <= 24'hd030c0;
             12'hd3d:  out <= 24'hd030d0;
             12'hd3e:  out <= 24'hd030e0;
             12'hd3f:  out <= 24'hd030f0;
             12'hd40:  out <= 24'hd04000;
             12'hd41:  out <= 24'hd04010;
             12'hd42:  out <= 24'hd04020;
             12'hd43:  out <= 24'hd04030;
             12'hd44:  out <= 24'hd04040;
             12'hd45:  out <= 24'hd04050;
             12'hd46:  out <= 24'hd04060;
             12'hd47:  out <= 24'hd04070;
             12'hd48:  out <= 24'hd04080;
             12'hd49:  out <= 24'hd04090;
             12'hd4a:  out <= 24'hd040a0;
             12'hd4b:  out <= 24'hd040b0;
             12'hd4c:  out <= 24'hd040c0;
             12'hd4d:  out <= 24'hd040d0;
             12'hd4e:  out <= 24'hd040e0;
             12'hd4f:  out <= 24'hd040f0;
             12'hd50:  out <= 24'hd05000;
             12'hd51:  out <= 24'hd05010;
             12'hd52:  out <= 24'hd05020;
             12'hd53:  out <= 24'hd05030;
             12'hd54:  out <= 24'hd05040;
             12'hd55:  out <= 24'hd05050;
             12'hd56:  out <= 24'hd05060;
             12'hd57:  out <= 24'hd05070;
             12'hd58:  out <= 24'hd05080;
             12'hd59:  out <= 24'hd05090;
             12'hd5a:  out <= 24'hd050a0;
             12'hd5b:  out <= 24'hd050b0;
             12'hd5c:  out <= 24'hd050c0;
             12'hd5d:  out <= 24'hd050d0;
             12'hd5e:  out <= 24'hd050e0;
             12'hd5f:  out <= 24'hd050f0;
             12'hd60:  out <= 24'hd06000;
             12'hd61:  out <= 24'hd06010;
             12'hd62:  out <= 24'hd06020;
             12'hd63:  out <= 24'hd06030;
             12'hd64:  out <= 24'hd06040;
             12'hd65:  out <= 24'hd06050;
             12'hd66:  out <= 24'hd06060;
             12'hd67:  out <= 24'hd06070;
             12'hd68:  out <= 24'hd06080;
             12'hd69:  out <= 24'hd06090;
             12'hd6a:  out <= 24'hd060a0;
             12'hd6b:  out <= 24'hd060b0;
             12'hd6c:  out <= 24'hd060c0;
             12'hd6d:  out <= 24'hd060d0;
             12'hd6e:  out <= 24'hd060e0;
             12'hd6f:  out <= 24'hd060f0;
             12'hd70:  out <= 24'hd07000;
             12'hd71:  out <= 24'hd07010;
             12'hd72:  out <= 24'hd07020;
             12'hd73:  out <= 24'hd07030;
             12'hd74:  out <= 24'hd07040;
             12'hd75:  out <= 24'hd07050;
             12'hd76:  out <= 24'hd07060;
             12'hd77:  out <= 24'hd07070;
             12'hd78:  out <= 24'hd07080;
             12'hd79:  out <= 24'hd07090;
             12'hd7a:  out <= 24'hd070a0;
             12'hd7b:  out <= 24'hd070b0;
             12'hd7c:  out <= 24'hd070c0;
             12'hd7d:  out <= 24'hd070d0;
             12'hd7e:  out <= 24'hd070e0;
             12'hd7f:  out <= 24'hd070f0;
             12'hd80:  out <= 24'hd08000;
             12'hd81:  out <= 24'hd08010;
             12'hd82:  out <= 24'hd08020;
             12'hd83:  out <= 24'hd08030;
             12'hd84:  out <= 24'hd08040;
             12'hd85:  out <= 24'hd08050;
             12'hd86:  out <= 24'hd08060;
             12'hd87:  out <= 24'hd08070;
             12'hd88:  out <= 24'hd08080;
             12'hd89:  out <= 24'hd08090;
             12'hd8a:  out <= 24'hd080a0;
             12'hd8b:  out <= 24'hd080b0;
             12'hd8c:  out <= 24'hd080c0;
             12'hd8d:  out <= 24'hd080d0;
             12'hd8e:  out <= 24'hd080e0;
             12'hd8f:  out <= 24'hd080f0;
             12'hd90:  out <= 24'hd09000;
             12'hd91:  out <= 24'hd09010;
             12'hd92:  out <= 24'hd09020;
             12'hd93:  out <= 24'hd09030;
             12'hd94:  out <= 24'hd09040;
             12'hd95:  out <= 24'hd09050;
             12'hd96:  out <= 24'hd09060;
             12'hd97:  out <= 24'hd09070;
             12'hd98:  out <= 24'hd09080;
             12'hd99:  out <= 24'hd09090;
             12'hd9a:  out <= 24'hd090a0;
             12'hd9b:  out <= 24'hd090b0;
             12'hd9c:  out <= 24'hd090c0;
             12'hd9d:  out <= 24'hd090d0;
             12'hd9e:  out <= 24'hd090e0;
             12'hd9f:  out <= 24'hd090f0;
             12'hda0:  out <= 24'hd0a000;
             12'hda1:  out <= 24'hd0a010;
             12'hda2:  out <= 24'hd0a020;
             12'hda3:  out <= 24'hd0a030;
             12'hda4:  out <= 24'hd0a040;
             12'hda5:  out <= 24'hd0a050;
             12'hda6:  out <= 24'hd0a060;
             12'hda7:  out <= 24'hd0a070;
             12'hda8:  out <= 24'hd0a080;
             12'hda9:  out <= 24'hd0a090;
             12'hdaa:  out <= 24'hd0a0a0;
             12'hdab:  out <= 24'hd0a0b0;
             12'hdac:  out <= 24'hd0a0c0;
             12'hdad:  out <= 24'hd0a0d0;
             12'hdae:  out <= 24'hd0a0e0;
             12'hdaf:  out <= 24'hd0a0f0;
             12'hdb0:  out <= 24'hd0b000;
             12'hdb1:  out <= 24'hd0b010;
             12'hdb2:  out <= 24'hd0b020;
             12'hdb3:  out <= 24'hd0b030;
             12'hdb4:  out <= 24'hd0b040;
             12'hdb5:  out <= 24'hd0b050;
             12'hdb6:  out <= 24'hd0b060;
             12'hdb7:  out <= 24'hd0b070;
             12'hdb8:  out <= 24'hd0b080;
             12'hdb9:  out <= 24'hd0b090;
             12'hdba:  out <= 24'hd0b0a0;
             12'hdbb:  out <= 24'hd0b0b0;
             12'hdbc:  out <= 24'hd0b0c0;
             12'hdbd:  out <= 24'hd0b0d0;
             12'hdbe:  out <= 24'hd0b0e0;
             12'hdbf:  out <= 24'hd0b0f0;
             12'hdc0:  out <= 24'hd0c000;
             12'hdc1:  out <= 24'hd0c010;
             12'hdc2:  out <= 24'hd0c020;
             12'hdc3:  out <= 24'hd0c030;
             12'hdc4:  out <= 24'hd0c040;
             12'hdc5:  out <= 24'hd0c050;
             12'hdc6:  out <= 24'hd0c060;
             12'hdc7:  out <= 24'hd0c070;
             12'hdc8:  out <= 24'hd0c080;
             12'hdc9:  out <= 24'hd0c090;
             12'hdca:  out <= 24'hd0c0a0;
             12'hdcb:  out <= 24'hd0c0b0;
             12'hdcc:  out <= 24'hd0c0c0;
             12'hdcd:  out <= 24'hd0c0d0;
             12'hdce:  out <= 24'hd0c0e0;
             12'hdcf:  out <= 24'hd0c0f0;
             12'hdd0:  out <= 24'hd0d000;
             12'hdd1:  out <= 24'hd0d010;
             12'hdd2:  out <= 24'hd0d020;
             12'hdd3:  out <= 24'hd0d030;
             12'hdd4:  out <= 24'hd0d040;
             12'hdd5:  out <= 24'hd0d050;
             12'hdd6:  out <= 24'hd0d060;
             12'hdd7:  out <= 24'hd0d070;
             12'hdd8:  out <= 24'hd0d080;
             12'hdd9:  out <= 24'hd0d090;
             12'hdda:  out <= 24'hd0d0a0;
             12'hddb:  out <= 24'hd0d0b0;
             12'hddc:  out <= 24'hd0d0c0;
             12'hddd:  out <= 24'hd0d0d0;
             12'hdde:  out <= 24'hd0d0e0;
             12'hddf:  out <= 24'hd0d0f0;
             12'hde0:  out <= 24'hd0e000;
             12'hde1:  out <= 24'hd0e010;
             12'hde2:  out <= 24'hd0e020;
             12'hde3:  out <= 24'hd0e030;
             12'hde4:  out <= 24'hd0e040;
             12'hde5:  out <= 24'hd0e050;
             12'hde6:  out <= 24'hd0e060;
             12'hde7:  out <= 24'hd0e070;
             12'hde8:  out <= 24'hd0e080;
             12'hde9:  out <= 24'hd0e090;
             12'hdea:  out <= 24'hd0e0a0;
             12'hdeb:  out <= 24'hd0e0b0;
             12'hdec:  out <= 24'hd0e0c0;
             12'hded:  out <= 24'hd0e0d0;
             12'hdee:  out <= 24'hd0e0e0;
             12'hdef:  out <= 24'hd0e0f0;
             12'hdf0:  out <= 24'hd0f000;
             12'hdf1:  out <= 24'hd0f010;
             12'hdf2:  out <= 24'hd0f020;
             12'hdf3:  out <= 24'hd0f030;
             12'hdf4:  out <= 24'hd0f040;
             12'hdf5:  out <= 24'hd0f050;
             12'hdf6:  out <= 24'hd0f060;
             12'hdf7:  out <= 24'hd0f070;
             12'hdf8:  out <= 24'hd0f080;
             12'hdf9:  out <= 24'hd0f090;
             12'hdfa:  out <= 24'hd0f0a0;
             12'hdfb:  out <= 24'hd0f0b0;
             12'hdfc:  out <= 24'hd0f0c0;
             12'hdfd:  out <= 24'hd0f0d0;
             12'hdfe:  out <= 24'hd0f0e0;
             12'hdff:  out <= 24'hd0f0f0;
             12'he00:  out <= 24'he00000;
             12'he01:  out <= 24'he00010;
             12'he02:  out <= 24'he00020;
             12'he03:  out <= 24'he00030;
             12'he04:  out <= 24'he00040;
             12'he05:  out <= 24'he00050;
             12'he06:  out <= 24'he00060;
             12'he07:  out <= 24'he00070;
             12'he08:  out <= 24'he00080;
             12'he09:  out <= 24'he00090;
             12'he0a:  out <= 24'he000a0;
             12'he0b:  out <= 24'he000b0;
             12'he0c:  out <= 24'he000c0;
             12'he0d:  out <= 24'he000d0;
             12'he0e:  out <= 24'he000e0;
             12'he0f:  out <= 24'he000f0;
             12'he10:  out <= 24'he01000;
             12'he11:  out <= 24'he01010;
             12'he12:  out <= 24'he01020;
             12'he13:  out <= 24'he01030;
             12'he14:  out <= 24'he01040;
             12'he15:  out <= 24'he01050;
             12'he16:  out <= 24'he01060;
             12'he17:  out <= 24'he01070;
             12'he18:  out <= 24'he01080;
             12'he19:  out <= 24'he01090;
             12'he1a:  out <= 24'he010a0;
             12'he1b:  out <= 24'he010b0;
             12'he1c:  out <= 24'he010c0;
             12'he1d:  out <= 24'he010d0;
             12'he1e:  out <= 24'he010e0;
             12'he1f:  out <= 24'he010f0;
             12'he20:  out <= 24'he02000;
             12'he21:  out <= 24'he02010;
             12'he22:  out <= 24'he02020;
             12'he23:  out <= 24'he02030;
             12'he24:  out <= 24'he02040;
             12'he25:  out <= 24'he02050;
             12'he26:  out <= 24'he02060;
             12'he27:  out <= 24'he02070;
             12'he28:  out <= 24'he02080;
             12'he29:  out <= 24'he02090;
             12'he2a:  out <= 24'he020a0;
             12'he2b:  out <= 24'he020b0;
             12'he2c:  out <= 24'he020c0;
             12'he2d:  out <= 24'he020d0;
             12'he2e:  out <= 24'he020e0;
             12'he2f:  out <= 24'he020f0;
             12'he30:  out <= 24'he03000;
             12'he31:  out <= 24'he03010;
             12'he32:  out <= 24'he03020;
             12'he33:  out <= 24'he03030;
             12'he34:  out <= 24'he03040;
             12'he35:  out <= 24'he03050;
             12'he36:  out <= 24'he03060;
             12'he37:  out <= 24'he03070;
             12'he38:  out <= 24'he03080;
             12'he39:  out <= 24'he03090;
             12'he3a:  out <= 24'he030a0;
             12'he3b:  out <= 24'he030b0;
             12'he3c:  out <= 24'he030c0;
             12'he3d:  out <= 24'he030d0;
             12'he3e:  out <= 24'he030e0;
             12'he3f:  out <= 24'he030f0;
             12'he40:  out <= 24'he04000;
             12'he41:  out <= 24'he04010;
             12'he42:  out <= 24'he04020;
             12'he43:  out <= 24'he04030;
             12'he44:  out <= 24'he04040;
             12'he45:  out <= 24'he04050;
             12'he46:  out <= 24'he04060;
             12'he47:  out <= 24'he04070;
             12'he48:  out <= 24'he04080;
             12'he49:  out <= 24'he04090;
             12'he4a:  out <= 24'he040a0;
             12'he4b:  out <= 24'he040b0;
             12'he4c:  out <= 24'he040c0;
             12'he4d:  out <= 24'he040d0;
             12'he4e:  out <= 24'he040e0;
             12'he4f:  out <= 24'he040f0;
             12'he50:  out <= 24'he05000;
             12'he51:  out <= 24'he05010;
             12'he52:  out <= 24'he05020;
             12'he53:  out <= 24'he05030;
             12'he54:  out <= 24'he05040;
             12'he55:  out <= 24'he05050;
             12'he56:  out <= 24'he05060;
             12'he57:  out <= 24'he05070;
             12'he58:  out <= 24'he05080;
             12'he59:  out <= 24'he05090;
             12'he5a:  out <= 24'he050a0;
             12'he5b:  out <= 24'he050b0;
             12'he5c:  out <= 24'he050c0;
             12'he5d:  out <= 24'he050d0;
             12'he5e:  out <= 24'he050e0;
             12'he5f:  out <= 24'he050f0;
             12'he60:  out <= 24'he06000;
             12'he61:  out <= 24'he06010;
             12'he62:  out <= 24'he06020;
             12'he63:  out <= 24'he06030;
             12'he64:  out <= 24'he06040;
             12'he65:  out <= 24'he06050;
             12'he66:  out <= 24'he06060;
             12'he67:  out <= 24'he06070;
             12'he68:  out <= 24'he06080;
             12'he69:  out <= 24'he06090;
             12'he6a:  out <= 24'he060a0;
             12'he6b:  out <= 24'he060b0;
             12'he6c:  out <= 24'he060c0;
             12'he6d:  out <= 24'he060d0;
             12'he6e:  out <= 24'he060e0;
             12'he6f:  out <= 24'he060f0;
             12'he70:  out <= 24'he07000;
             12'he71:  out <= 24'he07010;
             12'he72:  out <= 24'he07020;
             12'he73:  out <= 24'he07030;
             12'he74:  out <= 24'he07040;
             12'he75:  out <= 24'he07050;
             12'he76:  out <= 24'he07060;
             12'he77:  out <= 24'he07070;
             12'he78:  out <= 24'he07080;
             12'he79:  out <= 24'he07090;
             12'he7a:  out <= 24'he070a0;
             12'he7b:  out <= 24'he070b0;
             12'he7c:  out <= 24'he070c0;
             12'he7d:  out <= 24'he070d0;
             12'he7e:  out <= 24'he070e0;
             12'he7f:  out <= 24'he070f0;
             12'he80:  out <= 24'he08000;
             12'he81:  out <= 24'he08010;
             12'he82:  out <= 24'he08020;
             12'he83:  out <= 24'he08030;
             12'he84:  out <= 24'he08040;
             12'he85:  out <= 24'he08050;
             12'he86:  out <= 24'he08060;
             12'he87:  out <= 24'he08070;
             12'he88:  out <= 24'he08080;
             12'he89:  out <= 24'he08090;
             12'he8a:  out <= 24'he080a0;
             12'he8b:  out <= 24'he080b0;
             12'he8c:  out <= 24'he080c0;
             12'he8d:  out <= 24'he080d0;
             12'he8e:  out <= 24'he080e0;
             12'he8f:  out <= 24'he080f0;
             12'he90:  out <= 24'he09000;
             12'he91:  out <= 24'he09010;
             12'he92:  out <= 24'he09020;
             12'he93:  out <= 24'he09030;
             12'he94:  out <= 24'he09040;
             12'he95:  out <= 24'he09050;
             12'he96:  out <= 24'he09060;
             12'he97:  out <= 24'he09070;
             12'he98:  out <= 24'he09080;
             12'he99:  out <= 24'he09090;
             12'he9a:  out <= 24'he090a0;
             12'he9b:  out <= 24'he090b0;
             12'he9c:  out <= 24'he090c0;
             12'he9d:  out <= 24'he090d0;
             12'he9e:  out <= 24'he090e0;
             12'he9f:  out <= 24'he090f0;
             12'hea0:  out <= 24'he0a000;
             12'hea1:  out <= 24'he0a010;
             12'hea2:  out <= 24'he0a020;
             12'hea3:  out <= 24'he0a030;
             12'hea4:  out <= 24'he0a040;
             12'hea5:  out <= 24'he0a050;
             12'hea6:  out <= 24'he0a060;
             12'hea7:  out <= 24'he0a070;
             12'hea8:  out <= 24'he0a080;
             12'hea9:  out <= 24'he0a090;
             12'heaa:  out <= 24'he0a0a0;
             12'heab:  out <= 24'he0a0b0;
             12'heac:  out <= 24'he0a0c0;
             12'head:  out <= 24'he0a0d0;
             12'heae:  out <= 24'he0a0e0;
             12'heaf:  out <= 24'he0a0f0;
             12'heb0:  out <= 24'he0b000;
             12'heb1:  out <= 24'he0b010;
             12'heb2:  out <= 24'he0b020;
             12'heb3:  out <= 24'he0b030;
             12'heb4:  out <= 24'he0b040;
             12'heb5:  out <= 24'he0b050;
             12'heb6:  out <= 24'he0b060;
             12'heb7:  out <= 24'he0b070;
             12'heb8:  out <= 24'he0b080;
             12'heb9:  out <= 24'he0b090;
             12'heba:  out <= 24'he0b0a0;
             12'hebb:  out <= 24'he0b0b0;
             12'hebc:  out <= 24'he0b0c0;
             12'hebd:  out <= 24'he0b0d0;
             12'hebe:  out <= 24'he0b0e0;
             12'hebf:  out <= 24'he0b0f0;
             12'hec0:  out <= 24'he0c000;
             12'hec1:  out <= 24'he0c010;
             12'hec2:  out <= 24'he0c020;
             12'hec3:  out <= 24'he0c030;
             12'hec4:  out <= 24'he0c040;
             12'hec5:  out <= 24'he0c050;
             12'hec6:  out <= 24'he0c060;
             12'hec7:  out <= 24'he0c070;
             12'hec8:  out <= 24'he0c080;
             12'hec9:  out <= 24'he0c090;
             12'heca:  out <= 24'he0c0a0;
             12'hecb:  out <= 24'he0c0b0;
             12'hecc:  out <= 24'he0c0c0;
             12'hecd:  out <= 24'he0c0d0;
             12'hece:  out <= 24'he0c0e0;
             12'hecf:  out <= 24'he0c0f0;
             12'hed0:  out <= 24'he0d000;
             12'hed1:  out <= 24'he0d010;
             12'hed2:  out <= 24'he0d020;
             12'hed3:  out <= 24'he0d030;
             12'hed4:  out <= 24'he0d040;
             12'hed5:  out <= 24'he0d050;
             12'hed6:  out <= 24'he0d060;
             12'hed7:  out <= 24'he0d070;
             12'hed8:  out <= 24'he0d080;
             12'hed9:  out <= 24'he0d090;
             12'heda:  out <= 24'he0d0a0;
             12'hedb:  out <= 24'he0d0b0;
             12'hedc:  out <= 24'he0d0c0;
             12'hedd:  out <= 24'he0d0d0;
             12'hede:  out <= 24'he0d0e0;
             12'hedf:  out <= 24'he0d0f0;
             12'hee0:  out <= 24'he0e000;
             12'hee1:  out <= 24'he0e010;
             12'hee2:  out <= 24'he0e020;
             12'hee3:  out <= 24'he0e030;
             12'hee4:  out <= 24'he0e040;
             12'hee5:  out <= 24'he0e050;
             12'hee6:  out <= 24'he0e060;
             12'hee7:  out <= 24'he0e070;
             12'hee8:  out <= 24'he0e080;
             12'hee9:  out <= 24'he0e090;
             12'heea:  out <= 24'he0e0a0;
             12'heeb:  out <= 24'he0e0b0;
             12'heec:  out <= 24'he0e0c0;
             12'heed:  out <= 24'he0e0d0;
             12'heee:  out <= 24'he0e0e0;
             12'heef:  out <= 24'he0e0f0;
             12'hef0:  out <= 24'he0f000;
             12'hef1:  out <= 24'he0f010;
             12'hef2:  out <= 24'he0f020;
             12'hef3:  out <= 24'he0f030;
             12'hef4:  out <= 24'he0f040;
             12'hef5:  out <= 24'he0f050;
             12'hef6:  out <= 24'he0f060;
             12'hef7:  out <= 24'he0f070;
             12'hef8:  out <= 24'he0f080;
             12'hef9:  out <= 24'he0f090;
             12'hefa:  out <= 24'he0f0a0;
             12'hefb:  out <= 24'he0f0b0;
             12'hefc:  out <= 24'he0f0c0;
             12'hefd:  out <= 24'he0f0d0;
             12'hefe:  out <= 24'he0f0e0;
             12'heff:  out <= 24'he0f0f0;
             12'hf00:  out <= 24'hf00000;
             12'hf01:  out <= 24'hf00010;
             12'hf02:  out <= 24'hf00020;
             12'hf03:  out <= 24'hf00030;
             12'hf04:  out <= 24'hf00040;
             12'hf05:  out <= 24'hf00050;
             12'hf06:  out <= 24'hf00060;
             12'hf07:  out <= 24'hf00070;
             12'hf08:  out <= 24'hf00080;
             12'hf09:  out <= 24'hf00090;
             12'hf0a:  out <= 24'hf000a0;
             12'hf0b:  out <= 24'hf000b0;
             12'hf0c:  out <= 24'hf000c0;
             12'hf0d:  out <= 24'hf000d0;
             12'hf0e:  out <= 24'hf000e0;
             12'hf0f:  out <= 24'hf000f0;
             12'hf10:  out <= 24'hf01000;
             12'hf11:  out <= 24'hf01010;
             12'hf12:  out <= 24'hf01020;
             12'hf13:  out <= 24'hf01030;
             12'hf14:  out <= 24'hf01040;
             12'hf15:  out <= 24'hf01050;
             12'hf16:  out <= 24'hf01060;
             12'hf17:  out <= 24'hf01070;
             12'hf18:  out <= 24'hf01080;
             12'hf19:  out <= 24'hf01090;
             12'hf1a:  out <= 24'hf010a0;
             12'hf1b:  out <= 24'hf010b0;
             12'hf1c:  out <= 24'hf010c0;
             12'hf1d:  out <= 24'hf010d0;
             12'hf1e:  out <= 24'hf010e0;
             12'hf1f:  out <= 24'hf010f0;
             12'hf20:  out <= 24'hf02000;
             12'hf21:  out <= 24'hf02010;
             12'hf22:  out <= 24'hf02020;
             12'hf23:  out <= 24'hf02030;
             12'hf24:  out <= 24'hf02040;
             12'hf25:  out <= 24'hf02050;
             12'hf26:  out <= 24'hf02060;
             12'hf27:  out <= 24'hf02070;
             12'hf28:  out <= 24'hf02080;
             12'hf29:  out <= 24'hf02090;
             12'hf2a:  out <= 24'hf020a0;
             12'hf2b:  out <= 24'hf020b0;
             12'hf2c:  out <= 24'hf020c0;
             12'hf2d:  out <= 24'hf020d0;
             12'hf2e:  out <= 24'hf020e0;
             12'hf2f:  out <= 24'hf020f0;
             12'hf30:  out <= 24'hf03000;
             12'hf31:  out <= 24'hf03010;
             12'hf32:  out <= 24'hf03020;
             12'hf33:  out <= 24'hf03030;
             12'hf34:  out <= 24'hf03040;
             12'hf35:  out <= 24'hf03050;
             12'hf36:  out <= 24'hf03060;
             12'hf37:  out <= 24'hf03070;
             12'hf38:  out <= 24'hf03080;
             12'hf39:  out <= 24'hf03090;
             12'hf3a:  out <= 24'hf030a0;
             12'hf3b:  out <= 24'hf030b0;
             12'hf3c:  out <= 24'hf030c0;
             12'hf3d:  out <= 24'hf030d0;
             12'hf3e:  out <= 24'hf030e0;
             12'hf3f:  out <= 24'hf030f0;
             12'hf40:  out <= 24'hf04000;
             12'hf41:  out <= 24'hf04010;
             12'hf42:  out <= 24'hf04020;
             12'hf43:  out <= 24'hf04030;
             12'hf44:  out <= 24'hf04040;
             12'hf45:  out <= 24'hf04050;
             12'hf46:  out <= 24'hf04060;
             12'hf47:  out <= 24'hf04070;
             12'hf48:  out <= 24'hf04080;
             12'hf49:  out <= 24'hf04090;
             12'hf4a:  out <= 24'hf040a0;
             12'hf4b:  out <= 24'hf040b0;
             12'hf4c:  out <= 24'hf040c0;
             12'hf4d:  out <= 24'hf040d0;
             12'hf4e:  out <= 24'hf040e0;
             12'hf4f:  out <= 24'hf040f0;
             12'hf50:  out <= 24'hf05000;
             12'hf51:  out <= 24'hf05010;
             12'hf52:  out <= 24'hf05020;
             12'hf53:  out <= 24'hf05030;
             12'hf54:  out <= 24'hf05040;
             12'hf55:  out <= 24'hf05050;
             12'hf56:  out <= 24'hf05060;
             12'hf57:  out <= 24'hf05070;
             12'hf58:  out <= 24'hf05080;
             12'hf59:  out <= 24'hf05090;
             12'hf5a:  out <= 24'hf050a0;
             12'hf5b:  out <= 24'hf050b0;
             12'hf5c:  out <= 24'hf050c0;
             12'hf5d:  out <= 24'hf050d0;
             12'hf5e:  out <= 24'hf050e0;
             12'hf5f:  out <= 24'hf050f0;
             12'hf60:  out <= 24'hf06000;
             12'hf61:  out <= 24'hf06010;
             12'hf62:  out <= 24'hf06020;
             12'hf63:  out <= 24'hf06030;
             12'hf64:  out <= 24'hf06040;
             12'hf65:  out <= 24'hf06050;
             12'hf66:  out <= 24'hf06060;
             12'hf67:  out <= 24'hf06070;
             12'hf68:  out <= 24'hf06080;
             12'hf69:  out <= 24'hf06090;
             12'hf6a:  out <= 24'hf060a0;
             12'hf6b:  out <= 24'hf060b0;
             12'hf6c:  out <= 24'hf060c0;
             12'hf6d:  out <= 24'hf060d0;
             12'hf6e:  out <= 24'hf060e0;
             12'hf6f:  out <= 24'hf060f0;
             12'hf70:  out <= 24'hf07000;
             12'hf71:  out <= 24'hf07010;
             12'hf72:  out <= 24'hf07020;
             12'hf73:  out <= 24'hf07030;
             12'hf74:  out <= 24'hf07040;
             12'hf75:  out <= 24'hf07050;
             12'hf76:  out <= 24'hf07060;
             12'hf77:  out <= 24'hf07070;
             12'hf78:  out <= 24'hf07080;
             12'hf79:  out <= 24'hf07090;
             12'hf7a:  out <= 24'hf070a0;
             12'hf7b:  out <= 24'hf070b0;
             12'hf7c:  out <= 24'hf070c0;
             12'hf7d:  out <= 24'hf070d0;
             12'hf7e:  out <= 24'hf070e0;
             12'hf7f:  out <= 24'hf070f0;
             12'hf80:  out <= 24'hf08000;
             12'hf81:  out <= 24'hf08010;
             12'hf82:  out <= 24'hf08020;
             12'hf83:  out <= 24'hf08030;
             12'hf84:  out <= 24'hf08040;
             12'hf85:  out <= 24'hf08050;
             12'hf86:  out <= 24'hf08060;
             12'hf87:  out <= 24'hf08070;
             12'hf88:  out <= 24'hf08080;
             12'hf89:  out <= 24'hf08090;
             12'hf8a:  out <= 24'hf080a0;
             12'hf8b:  out <= 24'hf080b0;
             12'hf8c:  out <= 24'hf080c0;
             12'hf8d:  out <= 24'hf080d0;
             12'hf8e:  out <= 24'hf080e0;
             12'hf8f:  out <= 24'hf080f0;
             12'hf90:  out <= 24'hf09000;
             12'hf91:  out <= 24'hf09010;
             12'hf92:  out <= 24'hf09020;
             12'hf93:  out <= 24'hf09030;
             12'hf94:  out <= 24'hf09040;
             12'hf95:  out <= 24'hf09050;
             12'hf96:  out <= 24'hf09060;
             12'hf97:  out <= 24'hf09070;
             12'hf98:  out <= 24'hf09080;
             12'hf99:  out <= 24'hf09090;
             12'hf9a:  out <= 24'hf090a0;
             12'hf9b:  out <= 24'hf090b0;
             12'hf9c:  out <= 24'hf090c0;
             12'hf9d:  out <= 24'hf090d0;
             12'hf9e:  out <= 24'hf090e0;
             12'hf9f:  out <= 24'hf090f0;
             12'hfa0:  out <= 24'hf0a000;
             12'hfa1:  out <= 24'hf0a010;
             12'hfa2:  out <= 24'hf0a020;
             12'hfa3:  out <= 24'hf0a030;
             12'hfa4:  out <= 24'hf0a040;
             12'hfa5:  out <= 24'hf0a050;
             12'hfa6:  out <= 24'hf0a060;
             12'hfa7:  out <= 24'hf0a070;
             12'hfa8:  out <= 24'hf0a080;
             12'hfa9:  out <= 24'hf0a090;
             12'hfaa:  out <= 24'hf0a0a0;
             12'hfab:  out <= 24'hf0a0b0;
             12'hfac:  out <= 24'hf0a0c0;
             12'hfad:  out <= 24'hf0a0d0;
             12'hfae:  out <= 24'hf0a0e0;
             12'hfaf:  out <= 24'hf0a0f0;
             12'hfb0:  out <= 24'hf0b000;
             12'hfb1:  out <= 24'hf0b010;
             12'hfb2:  out <= 24'hf0b020;
             12'hfb3:  out <= 24'hf0b030;
             12'hfb4:  out <= 24'hf0b040;
             12'hfb5:  out <= 24'hf0b050;
             12'hfb6:  out <= 24'hf0b060;
             12'hfb7:  out <= 24'hf0b070;
             12'hfb8:  out <= 24'hf0b080;
             12'hfb9:  out <= 24'hf0b090;
             12'hfba:  out <= 24'hf0b0a0;
             12'hfbb:  out <= 24'hf0b0b0;
             12'hfbc:  out <= 24'hf0b0c0;
             12'hfbd:  out <= 24'hf0b0d0;
             12'hfbe:  out <= 24'hf0b0e0;
             12'hfbf:  out <= 24'hf0b0f0;
             12'hfc0:  out <= 24'hf0c000;
             12'hfc1:  out <= 24'hf0c010;
             12'hfc2:  out <= 24'hf0c020;
             12'hfc3:  out <= 24'hf0c030;
             12'hfc4:  out <= 24'hf0c040;
             12'hfc5:  out <= 24'hf0c050;
             12'hfc6:  out <= 24'hf0c060;
             12'hfc7:  out <= 24'hf0c070;
             12'hfc8:  out <= 24'hf0c080;
             12'hfc9:  out <= 24'hf0c090;
             12'hfca:  out <= 24'hf0c0a0;
             12'hfcb:  out <= 24'hf0c0b0;
             12'hfcc:  out <= 24'hf0c0c0;
             12'hfcd:  out <= 24'hf0c0d0;
             12'hfce:  out <= 24'hf0c0e0;
             12'hfcf:  out <= 24'hf0c0f0;
             12'hfd0:  out <= 24'hf0d000;
             12'hfd1:  out <= 24'hf0d010;
             12'hfd2:  out <= 24'hf0d020;
             12'hfd3:  out <= 24'hf0d030;
             12'hfd4:  out <= 24'hf0d040;
             12'hfd5:  out <= 24'hf0d050;
             12'hfd6:  out <= 24'hf0d060;
             12'hfd7:  out <= 24'hf0d070;
             12'hfd8:  out <= 24'hf0d080;
             12'hfd9:  out <= 24'hf0d090;
             12'hfda:  out <= 24'hf0d0a0;
             12'hfdb:  out <= 24'hf0d0b0;
             12'hfdc:  out <= 24'hf0d0c0;
             12'hfdd:  out <= 24'hf0d0d0;
             12'hfde:  out <= 24'hf0d0e0;
             12'hfdf:  out <= 24'hf0d0f0;
             12'hfe0:  out <= 24'hf0e000;
             12'hfe1:  out <= 24'hf0e010;
             12'hfe2:  out <= 24'hf0e020;
             12'hfe3:  out <= 24'hf0e030;
             12'hfe4:  out <= 24'hf0e040;
             12'hfe5:  out <= 24'hf0e050;
             12'hfe6:  out <= 24'hf0e060;
             12'hfe7:  out <= 24'hf0e070;
             12'hfe8:  out <= 24'hf0e080;
             12'hfe9:  out <= 24'hf0e090;
             12'hfea:  out <= 24'hf0e0a0;
             12'hfeb:  out <= 24'hf0e0b0;
             12'hfec:  out <= 24'hf0e0c0;
             12'hfed:  out <= 24'hf0e0d0;
             12'hfee:  out <= 24'hf0e0e0;
             12'hfef:  out <= 24'hf0e0f0;
             12'hff0:  out <= 24'hf0f000;
             12'hff1:  out <= 24'hf0f010;
             12'hff2:  out <= 24'hf0f020;
             12'hff3:  out <= 24'hf0f030;
             12'hff4:  out <= 24'hf0f040;
             12'hff5:  out <= 24'hf0f050;
             12'hff6:  out <= 24'hf0f060;
             12'hff7:  out <= 24'hf0f070;
             12'hff8:  out <= 24'hf0f080;
             12'hff9:  out <= 24'hf0f090;
             12'hffa:  out <= 24'hf0f0a0;
             12'hffb:  out <= 24'hf0f0b0;
             12'hffc:  out <= 24'hf0f0c0;
             12'hffd:  out <= 24'hf0f0d0;
             12'hffe:  out <= 24'hf0f0e0;
             12'hfff:  out <= 24'hf0f0f0;
        endcase
    end

endmodule