//-------------------------------------------------------------------------
//      lab8.sv                                                          --
//      Christine Chen                                                   --
//      Fall 2014                                                        --
//                                                                       --
//      Modified by Po-Han Huang                                         --
//      10/06/2017                                                       --
//                                                                       --
//      Fall 2017 Distribution                                           --
//                                                                       --
//      For use with ECE 385 Lab 8                                       --
//      UIUC ECE Department                                              --
//-------------------------------------------------------------------------


module top_level( 
            input               CLOCK_50,
            input        [3:0]  KEY,          //bit 0 is set up as Reset
            output logic [6:0]  HEX0, HEX1, HEX2, HEX3, HEX4, HEX5, HEX6, HEX7, // output to HEX displayer
            // VGA Interface 
            output logic [7:0]  VGA_R,        //VGA Red
                                VGA_G,        //VGA Green
                                VGA_B,        //VGA Blue
            output logic        VGA_CLK,      //VGA Clock
                                VGA_SYNC_N,   //VGA Sync signal
                                VGA_BLANK_N,  //VGA Blank signal
                                VGA_VS,       //VGA virtical sync signal
                                VGA_HS,       //VGA horizontal sync signal
            // CY7C67200 Interface
            inout  wire  [15:0] OTG_DATA,     //CY7C67200 Data bus 16 Bits
            output logic [1:0]  OTG_ADDR,     //CY7C67200 Address 2 Bits
            output logic        OTG_CS_N,     //CY7C67200 Chip Select
                                OTG_RD_N,     //CY7C67200 Write
                                OTG_WR_N,     //CY7C67200 Read
                                OTG_RST_N,    //CY7C67200 Reset
            input               OTG_INT,      //CY7C67200 Interrupt
            // SDRAM Interface for Nios II Software
            output logic [12:0] DRAM_ADDR,    //SDRAM Address 13 Bits
            inout  wire  [31:0] DRAM_DQ,      //SDRAM Data 32 Bits
            output logic [1:0]  DRAM_BA,      //SDRAM Bank Address 2 Bits
            output logic [3:0]  DRAM_DQM,     //SDRAM Data Mast 4 Bits
            output logic        DRAM_RAS_N,   //SDRAM Row Address Strobe
                                DRAM_CAS_N,   //SDRAM Column Address Strobe
                                DRAM_CKE,     //SDRAM Clock Enable
                                DRAM_WE_N,    //SDRAM Write Enable
                                DRAM_CS_N,    //SDRAM Chip Select
                                DRAM_CLK      //SDRAM Clock
                    );
    
    logic Reset_h, Clk;
    logic[9:0] DrawX, DrawY;
    
    assign Clk = CLOCK_50;
    always_ff @ (posedge Clk) begin
        Reset_h <= ~(KEY[0]);        // The push buttons are active low
    end
    
    logic [1:0] hpi_addr;
    logic [15:0] hpi_data_in, hpi_data_out;
    logic hpi_r, hpi_w, hpi_cs, hpi_reset;
    
    // Interface between NIOS II and EZ-OTG chip
    hpi_io_intf hpi_io_inst(
        .Clk(Clk),
        .Reset(Reset_h),
        // signals connected to NIOS II
        .from_sw_address(hpi_addr),
        .from_sw_data_in(hpi_data_in),
        .from_sw_data_out(hpi_data_out),
        .from_sw_r(hpi_r),
        .from_sw_w(hpi_w),
        .from_sw_cs(hpi_cs),
        .from_sw_reset(hpi_reset),
        // signals connected to EZ-OTG chip
        .OTG_DATA(OTG_DATA),    
        .OTG_ADDR(OTG_ADDR),    
        .OTG_RD_N(OTG_RD_N),    
        .OTG_WR_N(OTG_WR_N),    
        .OTG_CS_N(OTG_CS_N),
        .OTG_RST_N(OTG_RST_N)
    );
    logic [7:0] keycode_0, keycode_1, keycode_2, keycode_3, keycode_4, keycode_5, keycode_6, keycode_7;
     // You need to make sure that the port names here match the ports in Qsys-generated codes.
     final_soc nios_system(
        .clk_clk(Clk),         
        .reset_reset_n(1'b1),    // Never reset NIOS
        .sdram_wire_addr(DRAM_ADDR), 
        .sdram_wire_ba(DRAM_BA),   
        .sdram_wire_cas_n(DRAM_CAS_N),
        .sdram_wire_cke(DRAM_CKE),  
        .sdram_wire_cs_n(DRAM_CS_N), 
        .sdram_wire_dq(DRAM_DQ),   
        .sdram_wire_dqm(DRAM_DQM),  
        .sdram_wire_ras_n(DRAM_RAS_N),
        .sdram_wire_we_n(DRAM_WE_N), 
        .sdram_clk_clk(DRAM_CLK),

        .keycode_0_export(keycode_0),                              
        .keycode_1_export(keycode_1),  
        .keycode_2_export(keycode_2),
        .keycode_3_export(keycode_3),
        .keycode_4_export(keycode_4),  
        .keycode_5_export(keycode_5),

        .otg_hpi_address_export(hpi_addr),
        .otg_hpi_data_in_port(hpi_data_in),
        .otg_hpi_data_out_port(hpi_data_out),
        .otg_hpi_cs_export(hpi_cs),
        .otg_hpi_r_export(hpi_r),
        .otg_hpi_w_export(hpi_w),
        .otg_hpi_reset_export(hpi_reset)
    );
    
    // Use PLL to generate the 25MHZ VGA_CLK.
    // You will have to generate it on your own in simulation.
    vga_clk vga_clk_instance(.inclk0(Clk), .c0(VGA_CLK));
    
    VGA_controller vga_controller_instance(
        .Clk(Clk),
        .Reset(Reset_h),
        .VGA_HS,
        .VGA_VS,
        .VGA_CLK,
        .VGA_BLANK_N,
        .VGA_SYNC_N,
        .DrawX,
        .DrawY
    );
    
    wire [3:0] 	command_p1, command_p2; //{up, down, left, right}
    keycode u_keycode(
        //ports
        .Clk       		( Clk       		),
        .keycode_0 		( keycode_0 		),
        .keycode_1 		( keycode_1 		),
        .keycode_2 		( keycode_2 		),
        .keycode_3 		( keycode_3 		),
        .keycode_4 		( keycode_4 		),
        .keycode_5 		( keycode_5 		),

        .command_p1   	( command_p1   		),
        .command_p2     ( command_p2        )
    );

    wire [9:0] 	Ship_X_Step;
    wire       	Ship_Y_Step;
    wire [7:0] 	Ship_Angle;
    wire        forward;
    ship_controller #(
        .Ship_Max_Velocity_Forward 		( 10'd01 		),
        .Ship_Angle_Default        		( 8'b00010000   ))
    u_ship_controller(
        //ports
        .Clk         		( Clk         		),
        .Reset       		( Reset_h       	),
        .Command     		( command_p1     	),
        .Ship_X_Step 		( Ship_X_Step 		),
        .Ship_Y_Step 		( Ship_Y_Step 		),
        .Ship_Angle  		( Ship_Angle  		),
        .forward            ( forward           )
    );

    wire is_ball1;
    Ship #(
        .Ball_X_Center 		( 10'd480 		),
        .Ball_Y_Center 		( 10'd360 		),
        .Ball_X_Min    		( 10'd0   		),
        .Ball_X_Max    		( 10'd639 		),
        .Ball_Y_Min    		( 10'd0   		),
        .Ball_Y_Max    		( 10'd479 		),
        .Ball_Size     		( 10'd4   		))
    Ship_1(
        //ports
        .Clk       		( Clk       		),
        .Reset     		( Reset_h     		),
        .frame_clk 		( VGA_VS     		),
        .DrawX     		( DrawX     		),
        .DrawY     		( DrawY     		),
        .Step_X    		( Ship_X_Step    	),
        .Step_Y    		( Ship_Y_Step    	),
        .Angle     		( Ship_Angle     	),
        .is_ball   		( is_ball1   		)
    );

    wire [9:0] 	Ship_X_Step2;
    wire       	Ship_Y_Step2;
    wire [7:0] 	Ship_Angle2;
    wire        forward2;
    ship_controller #(
        .Ship_Max_Velocity_Forward 		( 10'd01 		),
        .Ship_Angle_Default        		( 8'b00000001   ))
    u_ship_controller2(
        //ports
        .Clk         		( Clk         		),
        .Reset       		( Reset_h       	),
        .Command     		( command_p2     	),
        .Ship_X_Step 		( Ship_X_Step2 		),
        .Ship_Y_Step 		( Ship_Y_Step2 		),
        .Ship_Angle  		( Ship_Angle2  		),
        .forward            ( forward2          )
    );

    wire is_ball2;
    Ship #(
        .Ball_X_Center 		( 10'd160 		),
        .Ball_Y_Center 		( 10'd120 		),
        .Ball_X_Min    		( 10'd0   		),
        .Ball_X_Max    		( 10'd639 		),
        .Ball_Y_Min    		( 10'd0   		),
        .Ball_Y_Max    		( 10'd479 		),
        .Ball_Size     		( 10'd4   		))
    Ship_2(
        //ports
        .Clk       		( Clk       		),
        .Reset     		( Reset_h     		),
        .frame_clk 		( VGA_VS     		),
        .DrawX     		( DrawX     		),
        .DrawY     		( DrawY     		),
        .Step_X    		( Ship_X_Step2    	),
        .Step_Y    		( Ship_Y_Step2    	),
        .Angle     		( Ship_Angle2     	),
        .is_ball   		( is_ball2   		)
    );

    logic [19:0] read_address;
    logic [7:0] bg_data, code;
    bgROM bg(.read_address, .Clk, .data_Out(bg_data));



    color_mapper u_color_mapper(
        //ports
        .is_ball1 		( is_ball1 		),
        .is_ball2 		( is_ball2 		),
        .code            ( code          ),
        .DrawX   		( DrawX   		),
        .DrawY   		( DrawY   		),
        .VGA_R   		( VGA_R   		),
        .VGA_G   		( VGA_G   		),
        .VGA_B   		( VGA_B   		)
    );


    // Display keycode on hex display
    HexDriver hex_inst_0 (Ship_Angle[3:0], HEX0);
    HexDriver hex_inst_1 (Ship_Angle[7:4], HEX1);
    HexDriver hex_inst_2 (Ship_Angle2[3:0], HEX2);
    HexDriver hex_inst_3 (Ship_Angle2[7:4], HEX3);


    always_comb
    begin
        code = bg_data;
    end
endmodule
